//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1184, new_n1185, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G77), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n203), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n207), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(G58), .A2(G68), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n221), .A2(G50), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G20), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n207), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n219), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G222), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(KEYINPUT68), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(KEYINPUT68), .B2(new_n258), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n267), .C1(G77), .C2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(G226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n224), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n283), .A2(new_n286), .B1(G150), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n204), .A2(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n281), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n280), .B1(new_n270), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(G50), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n278), .B(new_n296), .C1(G179), .C2(new_n276), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n276), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n296), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n276), .A2(G200), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n298), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT69), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n286), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n283), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n281), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n293), .A2(G77), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n291), .B2(G77), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n267), .A2(new_n273), .A3(new_n210), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n255), .A2(G232), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(new_n265), .C1(new_n216), .C2(new_n257), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G41), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n225), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n325), .B1(new_n328), .B2(new_n244), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n272), .B(new_n321), .C1(new_n323), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G190), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(G169), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n330), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n320), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n309), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n272), .B1(G238), .B2(new_n274), .ZN(new_n341));
  OR2_X1    g0141(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G226), .A3(new_n252), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G232), .A2(G1698), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n328), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n267), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n341), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n341), .A2(new_n348), .A3(KEYINPUT73), .A4(new_n349), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n341), .B2(new_n348), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(G179), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n350), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT14), .B1(new_n358), .B2(G169), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n360), .B(new_n277), .C1(new_n356), .C2(new_n350), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n203), .A2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(new_n287), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n363), .B1(new_n285), .B2(new_n209), .C1(new_n364), .C2(new_n201), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n280), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT11), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT11), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n366), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT75), .ZN(new_n372));
  INV_X1    g0172(.A(new_n293), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT12), .B1(new_n373), .B2(new_n203), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n373), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(G68), .C2(new_n291), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n362), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n358), .A2(new_n379), .A3(G200), .ZN(new_n380));
  INV_X1    g0180(.A(new_n350), .ZN(new_n381));
  OAI21_X1  g0181(.A(G200), .B1(new_n381), .B2(new_n355), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT72), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n355), .A2(new_n300), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n354), .A2(KEYINPUT74), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n352), .A3(new_n353), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n378), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n263), .A2(new_n284), .A3(new_n264), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n284), .A4(new_n264), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT76), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G68), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n202), .A2(new_n203), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n220), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n287), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n281), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n203), .B1(new_n395), .B2(new_n396), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n408), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT77), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT77), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n405), .C1(new_n408), .C2(new_n404), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n342), .A2(G223), .A3(new_n252), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G226), .A2(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n328), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n267), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n269), .B1(new_n225), .B2(new_n324), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n273), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n325), .A2(G232), .A3(new_n271), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n332), .ZN(new_n425));
  AND2_X1   g0225(.A1(KEYINPUT80), .A2(G190), .ZN(new_n426));
  NOR2_X1   g0226(.A1(KEYINPUT80), .A2(G190), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n421), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n421), .B2(new_n422), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n419), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n283), .A2(new_n293), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n291), .B2(new_n283), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n413), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n413), .A2(new_n438), .A3(new_n433), .A4(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n413), .A2(new_n435), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n430), .A2(new_n431), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(KEYINPUT79), .A3(new_n337), .A4(new_n419), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n419), .B(new_n337), .C1(new_n430), .C2(new_n431), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n424), .A2(new_n277), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT18), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n413), .A2(new_n435), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n446), .A2(new_n447), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n443), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n440), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n373), .A2(new_n246), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n270), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n281), .A2(G116), .A3(new_n293), .A4(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n279), .A2(new_n224), .B1(G20), .B2(new_n246), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n284), .C1(G33), .C2(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT20), .B1(new_n458), .B2(new_n461), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n455), .B(new_n457), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G41), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n270), .B(G45), .C1(new_n466), .C2(KEYINPUT5), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n420), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n325), .B(G270), .C1(new_n467), .C2(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G264), .A2(G1698), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n326), .B2(new_n327), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(G257), .B2(new_n255), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n267), .B1(new_n265), .B2(G303), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n470), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n465), .A2(new_n337), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n464), .A3(G169), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT21), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n476), .A2(new_n464), .A3(new_n480), .A4(G169), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G257), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n257), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n265), .A2(new_n484), .B1(G33), .B2(G294), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n212), .B1(new_n263), .B2(new_n264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n255), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n325), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n325), .B(G264), .C1(new_n467), .C2(new_n468), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n470), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(G169), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n488), .A2(new_n490), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n337), .ZN(new_n493));
  AOI21_X1  g0293(.A(G20), .B1(new_n263), .B2(new_n264), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT22), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(G87), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n284), .B(G87), .C1(new_n326), .C2(new_n327), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT22), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OR3_X1    g0299(.A1(new_n284), .A2(KEYINPUT23), .A3(G107), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT87), .B1(new_n501), .B2(G20), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT23), .B1(new_n284), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n501), .A2(KEYINPUT87), .A3(G20), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT24), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n499), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n281), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n373), .A2(new_n244), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n512), .A2(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(KEYINPUT25), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n281), .A2(new_n293), .A3(new_n456), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n244), .C2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n493), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n499), .A2(new_n509), .A3(new_n506), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n509), .B1(new_n499), .B2(new_n506), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n280), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n492), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  OR3_X1    g0322(.A1(new_n488), .A2(new_n490), .A3(new_n300), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n476), .A2(G200), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n525), .B(new_n465), .C1(new_n428), .C2(new_n476), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n482), .A2(new_n517), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n342), .A2(G238), .A3(new_n252), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G244), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n328), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n501), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n267), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n270), .A2(new_n269), .A3(G45), .ZN(new_n533));
  INV_X1    g0333(.A(G45), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n212), .B1(new_n534), .B2(G1), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n325), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(KEYINPUT84), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT84), .B1(new_n532), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g0339(.A(G200), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n532), .A2(new_n536), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT84), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n537), .A3(G190), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n312), .A2(new_n293), .ZN(new_n545));
  NOR3_X1   g0345(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n284), .B1(new_n547), .B2(new_n346), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(KEYINPUT86), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n284), .C1(new_n547), .C2(new_n346), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n494), .A2(G68), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n547), .B1(new_n460), .B2(new_n285), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n545), .B1(new_n557), .B2(new_n280), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n515), .A2(new_n211), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n540), .A2(new_n544), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n277), .B1(new_n538), .B2(new_n539), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n543), .A2(new_n537), .A3(new_n337), .ZN(new_n563));
  INV_X1    g0363(.A(new_n545), .ZN(new_n564));
  INV_X1    g0364(.A(new_n515), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n312), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n555), .B1(new_n549), .B2(new_n551), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n566), .C1(new_n567), .C2(new_n281), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n527), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n210), .B1(new_n263), .B2(new_n264), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(KEYINPUT4), .A3(new_n255), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT81), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n255), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT81), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n572), .A2(new_n255), .A3(new_n578), .A4(KEYINPUT4), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n486), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n574), .A2(new_n577), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n267), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n325), .B(G257), .C1(new_n467), .C2(new_n468), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n470), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(KEYINPUT82), .A3(G200), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n244), .A2(KEYINPUT6), .A3(G97), .ZN(new_n588));
  XNOR2_X1  g0388(.A(G97), .B(G107), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n591), .A2(new_n284), .B1(new_n209), .B2(new_n364), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n244), .B1(new_n395), .B2(new_n396), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n280), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n293), .A2(G97), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n565), .B2(G97), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n584), .B1(new_n581), .B2(new_n267), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(G190), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT82), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n598), .B2(new_n332), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n587), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n337), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(new_n597), .C1(G169), .C2(new_n598), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n602), .A2(KEYINPUT83), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT83), .B1(new_n602), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n571), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR4_X1   g0407(.A1(new_n340), .A2(new_n392), .A3(new_n454), .A4(new_n607), .ZN(G372));
  NOR3_X1   g0408(.A1(new_n340), .A2(new_n392), .A3(new_n454), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT26), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n570), .A2(new_n610), .A3(new_n604), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n602), .A2(new_n604), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n559), .B1(new_n541), .B2(G200), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n544), .A2(new_n558), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n541), .A2(new_n277), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n563), .A2(new_n568), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n482), .A2(new_n517), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n614), .A2(new_n524), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n613), .A2(new_n622), .A3(new_n618), .ZN(new_n623));
  INV_X1    g0423(.A(new_n604), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT26), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n625), .A2(new_n611), .A3(new_n612), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n449), .A2(new_n453), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n339), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n377), .B2(new_n362), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n391), .A2(new_n440), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n307), .A2(new_n308), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n298), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n628), .A2(new_n636), .ZN(G369));
  INV_X1    g0437(.A(new_n482), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n270), .A2(new_n284), .A3(G13), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n465), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n482), .A2(new_n526), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n646), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n517), .A2(new_n524), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n644), .B1(new_n511), .B2(new_n516), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n517), .B2(new_n645), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n482), .A2(new_n644), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n517), .B2(new_n644), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(G399));
  NAND2_X1  g0461(.A1(new_n546), .A2(new_n246), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT89), .Z(new_n663));
  INV_X1    g0463(.A(new_n228), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n663), .A2(new_n270), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n223), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n665), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT28), .Z(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n627), .A2(new_n670), .A3(new_n645), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n622), .A2(new_n618), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n619), .B2(new_n604), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n624), .A2(new_n569), .A3(new_n561), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(KEYINPUT26), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n645), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT29), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n571), .B(new_n645), .C1(new_n605), .C2(new_n606), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT91), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n681), .A2(new_n488), .A3(new_n490), .A4(new_n337), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n598), .A3(new_n543), .A4(new_n537), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(KEYINPUT90), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n683), .B2(KEYINPUT90), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n492), .A2(new_n541), .A3(new_n337), .A4(new_n476), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n598), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n645), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n680), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n690), .B1(new_n689), .B2(new_n645), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n686), .A2(new_n688), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n683), .A2(KEYINPUT90), .A3(new_n684), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT91), .A3(new_n691), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n679), .A2(new_n693), .A3(new_n694), .A4(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n678), .B1(G330), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n669), .B1(new_n700), .B2(G1), .ZN(G364));
  INV_X1    g0501(.A(new_n665), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n284), .A2(G13), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n270), .B1(new_n703), .B2(G45), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n649), .A2(G330), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n651), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT92), .Z(new_n709));
  NOR2_X1   g0509(.A1(new_n664), .A2(new_n328), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G355), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G116), .B2(new_n228), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n664), .A2(new_n265), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n667), .B2(new_n534), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n250), .A2(G45), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT93), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n224), .B1(G20), .B2(new_n277), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n706), .B1(new_n717), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n720), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n649), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n284), .A2(new_n337), .A3(new_n332), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT95), .A3(new_n300), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT95), .B1(new_n727), .B2(new_n300), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n428), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n284), .A2(new_n337), .A3(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n300), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n202), .B1(new_n209), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT94), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n731), .A2(G68), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n737), .B2(new_n736), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n284), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n300), .A3(new_n332), .ZN(new_n741));
  INV_X1    g0541(.A(G159), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT32), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n732), .A2(new_n727), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n328), .B1(new_n746), .B2(G50), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G87), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n300), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n284), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n740), .A2(new_n300), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n753), .A2(G97), .B1(new_n755), .B2(G107), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n744), .A2(new_n747), .A3(new_n750), .A4(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n745), .B(KEYINPUT96), .Z(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT33), .B(G317), .Z(new_n760));
  OAI22_X1  g0560(.A1(new_n758), .A2(new_n759), .B1(new_n730), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n734), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G322), .ZN(new_n763));
  INV_X1    g0563(.A(new_n735), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G311), .B1(new_n755), .B2(G283), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n753), .A2(G294), .B1(new_n749), .B2(G303), .ZN(new_n766));
  INV_X1    g0566(.A(new_n741), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n265), .B1(new_n767), .B2(G329), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n763), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n739), .A2(new_n757), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n724), .B(new_n726), .C1(new_n721), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n709), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  NAND2_X1  g0573(.A1(new_n320), .A2(new_n644), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n631), .B1(new_n335), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n339), .A2(new_n644), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n627), .B2(new_n645), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n645), .C1(new_n623), .C2(new_n626), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n699), .A2(G330), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n706), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n721), .A2(new_n718), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n706), .B1(G77), .B2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n762), .A2(G143), .B1(G159), .B2(new_n764), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n745), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G150), .B2(new_n731), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n792));
  INV_X1    g0592(.A(G132), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n265), .B1(new_n741), .B2(new_n793), .C1(new_n201), .C2(new_n748), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n752), .A2(new_n202), .B1(new_n754), .B2(new_n203), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(KEYINPUT34), .B2(new_n791), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n746), .A2(G303), .B1(G116), .B2(new_n764), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n730), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT97), .Z(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n328), .B1(new_n741), .B2(new_n802), .C1(new_n752), .C2(new_n460), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n734), .A2(new_n804), .B1(new_n244), .B2(new_n748), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(G87), .C2(new_n755), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n787), .B1(new_n808), .B2(new_n721), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT98), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n719), .B2(new_n777), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n784), .A2(new_n811), .ZN(G384));
  INV_X1    g0612(.A(new_n591), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT35), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n226), .A2(new_n246), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n813), .B2(KEYINPUT35), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT36), .ZN(new_n820));
  OR3_X1    g0620(.A1(new_n223), .A2(new_n209), .A3(new_n401), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n201), .A2(G68), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n270), .B(G13), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n703), .A2(new_n270), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n378), .A2(new_n644), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n435), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n405), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n407), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n436), .B1(new_n831), .B2(new_n642), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n448), .A2(new_n831), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT37), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n642), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n450), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n836), .B(new_n436), .C1(new_n441), .C2(new_n448), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n834), .B1(KEYINPUT37), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT101), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n831), .A2(new_n642), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n454), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n454), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(KEYINPUT38), .B(new_n838), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(KEYINPUT102), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n843), .A2(new_n848), .A3(new_n844), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(KEYINPUT39), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n837), .B(KEYINPUT37), .Z(new_n851));
  AOI21_X1  g0651(.A(new_n836), .B1(new_n630), .B2(new_n440), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(new_n846), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n827), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n377), .A2(new_n644), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n378), .A2(new_n391), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n362), .A2(new_n377), .A3(new_n644), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT100), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n776), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n779), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n847), .A2(new_n849), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n629), .A2(new_n642), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n856), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n678), .A2(new_n609), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n636), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n870), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n697), .A2(new_n691), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n694), .A2(new_n679), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n858), .A2(new_n862), .A3(new_n859), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n862), .B1(new_n858), .B2(new_n859), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n777), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n847), .A2(new_n849), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n853), .B2(new_n846), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n880), .A2(new_n881), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n609), .A2(new_n875), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  INV_X1    g0686(.A(G330), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n825), .B1(new_n873), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT103), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n889), .A2(new_n890), .B1(new_n873), .B2(new_n888), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n824), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT104), .ZN(G367));
  NAND2_X1  g0694(.A1(new_n597), .A2(new_n644), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n614), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT105), .Z(new_n897));
  NAND2_X1  g0697(.A1(new_n624), .A2(new_n644), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n652), .A3(new_n657), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n604), .B1(new_n897), .B2(new_n517), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n900), .A2(KEYINPUT42), .B1(new_n901), .B2(new_n645), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(KEYINPUT42), .B2(new_n900), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n645), .B1(new_n558), .B2(new_n560), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n568), .A3(new_n563), .A4(new_n617), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n619), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n656), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n899), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n908), .B(new_n909), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n899), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n665), .B(KEYINPUT41), .Z(new_n916));
  INV_X1    g0716(.A(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n899), .A2(new_n660), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n899), .A2(new_n660), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT44), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(KEYINPUT107), .A3(new_n911), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n658), .B1(new_n655), .B2(new_n657), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(new_n651), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n700), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n921), .A2(new_n924), .A3(new_n933), .A4(new_n926), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n928), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n916), .B1(new_n935), .B2(new_n700), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n704), .B(KEYINPUT108), .Z(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n912), .B(new_n915), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n723), .B1(new_n240), .B2(new_n713), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n312), .A2(new_n664), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n762), .A2(G303), .B1(G283), .B2(new_n764), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n244), .B2(new_n752), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(G294), .B2(new_n731), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n749), .A2(KEYINPUT46), .A3(G116), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT46), .B1(new_n749), .B2(G116), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n754), .A2(new_n460), .ZN(new_n948));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n328), .B1(new_n741), .B2(new_n949), .ZN(new_n950));
  NOR4_X1   g0750(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n945), .B(new_n951), .C1(new_n802), .C2(new_n758), .ZN(new_n952));
  INV_X1    g0752(.A(G150), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n265), .B1(new_n789), .B2(new_n741), .C1(new_n734), .C2(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n202), .A2(new_n748), .B1(new_n754), .B2(new_n209), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n735), .A2(new_n201), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n752), .A2(new_n203), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(G143), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n958), .B1(new_n959), .B2(new_n758), .C1(new_n742), .C2(new_n730), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n952), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n705), .B(new_n942), .C1(new_n962), .C2(new_n721), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n906), .B2(new_n725), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n939), .A2(new_n964), .ZN(G387));
  NOR2_X1   g0765(.A1(new_n932), .A2(new_n702), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n700), .B2(new_n930), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n930), .A2(new_n938), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT109), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n328), .B(new_n948), .C1(G150), .C2(new_n767), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n748), .A2(new_n209), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n762), .B2(G50), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n746), .A2(G159), .B1(G68), .B2(new_n764), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n312), .A2(new_n753), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n283), .B2(new_n731), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT112), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n265), .B1(new_n767), .B2(G326), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n752), .A2(new_n799), .B1(new_n748), .B2(new_n804), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n762), .A2(G317), .B1(G303), .B2(new_n764), .ZN(new_n980));
  INV_X1    g0780(.A(G322), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n980), .B1(new_n802), .B2(new_n730), .C1(new_n758), .C2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT48), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT49), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n978), .B1(new_n246), .B2(new_n754), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n721), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n655), .A2(new_n725), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n714), .B1(new_n237), .B2(G45), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT111), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n663), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n282), .A2(KEYINPUT50), .A3(G50), .ZN(new_n995));
  AOI211_X1 g0795(.A(G45), .B(new_n995), .C1(G68), .C2(G77), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n663), .A2(new_n993), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT50), .B1(new_n282), .B2(G50), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n992), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n663), .A2(new_n710), .B1(new_n244), .B2(new_n664), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT110), .Z(new_n1002));
  AOI21_X1  g0802(.A(new_n723), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n991), .A2(new_n705), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n969), .B1(new_n990), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n967), .A2(new_n1005), .ZN(G393));
  NAND2_X1  g0806(.A1(new_n927), .A2(new_n911), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n921), .A2(new_n924), .A3(new_n656), .A4(new_n926), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n938), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n247), .A2(new_n714), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n722), .B1(new_n460), .B2(new_n228), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n706), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n265), .B1(new_n741), .B2(new_n959), .C1(new_n211), .C2(new_n754), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n753), .A2(G77), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n282), .B2(new_n735), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G68), .C2(new_n749), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n201), .B2(new_n730), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n953), .A2(new_n745), .B1(new_n734), .B2(new_n742), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT51), .Z(new_n1019));
  OAI22_X1  g0819(.A1(new_n802), .A2(new_n734), .B1(new_n745), .B2(new_n949), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT52), .Z(new_n1021));
  OAI22_X1  g0821(.A1(new_n735), .A2(new_n804), .B1(new_n752), .B2(new_n246), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n328), .B1(new_n741), .B2(new_n981), .C1(new_n244), .C2(new_n754), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G283), .C2(new_n749), .ZN(new_n1024));
  INV_X1    g0824(.A(G303), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n730), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1017), .A2(new_n1019), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n1012), .B1(new_n1028), .B2(new_n721), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n899), .B2(new_n725), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1009), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n935), .A2(new_n665), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n931), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1031), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G390));
  AND2_X1   g0836(.A1(new_n875), .A2(G330), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n609), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n871), .A2(new_n636), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n699), .A2(G330), .A3(new_n777), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n876), .A2(new_n877), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(new_n777), .A3(new_n864), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT115), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1040), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n866), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT114), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n864), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1037), .A2(new_n777), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1040), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n864), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n676), .A2(new_n775), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1057), .A2(new_n865), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1039), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n866), .A2(new_n864), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n827), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n850), .A2(new_n1063), .A3(new_n855), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n826), .B1(new_n853), .B2(new_n846), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1058), .B2(new_n1052), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1056), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1044), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1061), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1044), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n1060), .A3(new_n1067), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1070), .A2(new_n665), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n706), .B1(new_n283), .B2(new_n786), .ZN(new_n1076));
  INV_X1    g0876(.A(G128), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n745), .A2(new_n1077), .B1(new_n201), .B2(new_n754), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n328), .B1(new_n767), .B2(G125), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n793), .B2(new_n734), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(G159), .C2(new_n753), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n735), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n731), .B2(G137), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n748), .A2(new_n953), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT53), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1081), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n746), .A2(G283), .B1(G97), .B2(new_n764), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n730), .B2(new_n244), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n762), .A2(G116), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1093), .A2(new_n328), .A3(new_n750), .A4(new_n1014), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n754), .A2(new_n203), .B1(new_n741), .B2(new_n804), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT119), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1088), .A2(new_n1089), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1076), .B1(new_n1098), .B2(new_n721), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n850), .A2(new_n855), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n719), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n938), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT116), .A4(new_n937), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1075), .B(new_n1101), .C1(new_n1104), .C2(new_n1105), .ZN(G378));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n826), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n869), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n880), .A2(new_n881), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n887), .B1(new_n882), .B2(new_n879), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n309), .B(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n296), .A2(new_n835), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1110), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1109), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1110), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1116), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n870), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n937), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n706), .B1(G50), .B2(new_n786), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1117), .A2(new_n719), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n265), .A2(G41), .ZN(new_n1127));
  AOI211_X1 g0927(.A(G50), .B(new_n1127), .C1(new_n262), .C2(new_n466), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n244), .A2(new_n734), .B1(new_n745), .B2(new_n246), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n971), .B(new_n1129), .C1(G58), .C2(new_n755), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n799), .B2(new_n741), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n957), .B(new_n1131), .C1(new_n312), .C2(new_n764), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n460), .C2(new_n730), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT58), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1128), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n748), .A2(new_n1082), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT120), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n746), .A2(G125), .B1(G150), .B2(new_n753), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n1077), .B2(new_n734), .C1(new_n789), .C2(new_n735), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G132), .C2(new_n731), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT59), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1136), .B1(new_n742), .B2(new_n754), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1135), .B1(new_n1134), .B2(new_n1133), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1125), .B(new_n1126), .C1(new_n721), .C2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1124), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1120), .A2(new_n1123), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1039), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1074), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1109), .A2(new_n1118), .A3(KEYINPUT121), .A4(new_n1119), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT57), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1153), .A2(KEYINPUT57), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1147), .B1(new_n1155), .B2(new_n702), .ZN(G375));
  INV_X1    g0956(.A(new_n916), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1048), .A2(new_n1039), .A3(new_n1059), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1061), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n937), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1052), .A2(new_n718), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n706), .B1(G68), .B2(new_n786), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n762), .A2(G137), .B1(G50), .B2(new_n753), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n742), .B2(new_n748), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n265), .B1(new_n741), .B2(new_n1077), .C1(new_n202), .C2(new_n754), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n745), .A2(new_n793), .B1(new_n953), .B2(new_n735), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n730), .B2(new_n1082), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G283), .A2(new_n762), .B1(new_n746), .B2(G294), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n764), .A2(G107), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n265), .B1(new_n755), .B2(G77), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n974), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n741), .A2(new_n1025), .B1(new_n748), .B2(new_n460), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n731), .A2(G116), .B1(KEYINPUT122), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(KEYINPUT122), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1168), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1162), .B1(new_n1176), .B2(new_n721), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1160), .B1(new_n1161), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n1178), .ZN(G381));
  NAND3_X1  g0979(.A1(new_n939), .A2(new_n1035), .A3(new_n964), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n967), .A2(new_n772), .A3(new_n1005), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1181), .A2(G381), .A3(G384), .ZN(new_n1182));
  OR4_X1    g0982(.A1(G378), .A2(G375), .A3(new_n1180), .A4(new_n1182), .ZN(G407));
  NAND2_X1  g0983(.A1(new_n643), .A2(G213), .ZN(new_n1184));
  OR3_X1    g0984(.A1(G375), .A2(G378), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(G407), .A2(G213), .A3(new_n1185), .ZN(G409));
  OAI211_X1 g0986(.A(G378), .B(new_n1147), .C1(new_n1155), .C2(new_n702), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n916), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT123), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1151), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1189), .B2(new_n1151), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1146), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT124), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT124), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1149), .A2(new_n1196), .A3(new_n1152), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n938), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G378), .B1(new_n1193), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1184), .B1(new_n1188), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT127), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1060), .A2(new_n702), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT60), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1158), .A2(KEYINPUT125), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n1158), .B2(KEYINPUT125), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G384), .B(new_n1178), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1158), .A2(KEYINPUT125), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n1204), .A3(new_n1202), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G384), .B1(new_n1211), .B2(new_n1178), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n643), .A2(G213), .A3(G2897), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1201), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  OAI211_X1 g1016(.A(KEYINPUT127), .B(new_n1216), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1211), .A2(new_n1178), .ZN(new_n1218));
  INV_X1    g1018(.A(G384), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1207), .A3(new_n1214), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(KEYINPUT126), .A3(new_n1207), .A4(new_n1214), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1215), .A2(new_n1217), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT61), .B1(new_n1200), .B2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1187), .B1(new_n1227), .B2(G378), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT62), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1184), .A4(new_n1213), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1184), .B(new_n1213), .C1(new_n1188), .C2(new_n1199), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT62), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1226), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1180), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1035), .B1(new_n939), .B2(new_n964), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1181), .B(new_n1234), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(G390), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1181), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1180), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1233), .A2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1228), .A2(KEYINPUT63), .A3(new_n1184), .A4(new_n1213), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1231), .A2(new_n1244), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1238), .A2(new_n1180), .A3(new_n1239), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1239), .B1(new_n1238), .B2(new_n1180), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1226), .A2(new_n1243), .A3(new_n1245), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1249), .ZN(G405));
  INV_X1    g1050(.A(new_n1213), .ZN(new_n1251));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G375), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1187), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1241), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1251), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1241), .A2(new_n1256), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1213), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(G402));
endmodule


