

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U550 ( .A(n896), .Z(n518) );
  INV_X1 U551 ( .A(n743), .ZN(n764) );
  INV_X1 U552 ( .A(G2105), .ZN(n525) );
  BUF_X1 U553 ( .A(n892), .Z(n517) );
  NOR2_X1 U554 ( .A1(G2104), .A2(n525), .ZN(n892) );
  AND2_X1 U555 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U557 ( .A(n527), .B(n526), .ZN(n896) );
  NAND2_X1 U558 ( .A1(G40), .A2(G160), .ZN(n711) );
  AND2_X1 U559 ( .A1(n777), .A2(n519), .ZN(n778) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n710) );
  INV_X1 U561 ( .A(KEYINPUT17), .ZN(n526) );
  NOR2_X2 U562 ( .A1(n636), .A2(n544), .ZN(n652) );
  NOR2_X1 U563 ( .A1(n776), .A2(n775), .ZN(n519) );
  NOR2_X4 U564 ( .A1(n712), .A2(n711), .ZN(n743) );
  XNOR2_X1 U565 ( .A(KEYINPUT28), .B(n740), .ZN(n520) );
  AND2_X1 U566 ( .A1(n741), .A2(n520), .ZN(n521) );
  INV_X1 U567 ( .A(KEYINPUT26), .ZN(n724) );
  INV_X1 U568 ( .A(KEYINPUT30), .ZN(n752) );
  INV_X1 U569 ( .A(KEYINPUT94), .ZN(n713) );
  INV_X1 U570 ( .A(n715), .ZN(n799) );
  INV_X1 U571 ( .A(KEYINPUT73), .ZN(n594) );
  XNOR2_X1 U572 ( .A(n594), .B(KEYINPUT13), .ZN(n595) );
  NAND2_X1 U573 ( .A1(n896), .A2(G137), .ZN(n532) );
  XNOR2_X1 U574 ( .A(n596), .B(n595), .ZN(n600) );
  NOR2_X1 U575 ( .A1(G651), .A2(n636), .ZN(n657) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U577 ( .A1(n602), .A2(n601), .ZN(n1006) );
  NOR2_X1 U578 ( .A1(n531), .A2(n530), .ZN(G164) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U580 ( .A1(G114), .A2(n891), .ZN(n523) );
  NAND2_X1 U581 ( .A1(G126), .A2(n892), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U583 ( .A(KEYINPUT86), .B(n524), .ZN(n531) );
  AND2_X4 U584 ( .A1(n525), .A2(G2104), .ZN(n895) );
  NAND2_X1 U585 ( .A1(G102), .A2(n895), .ZN(n529) );
  NAND2_X1 U586 ( .A1(G138), .A2(n518), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n892), .A2(G125), .ZN(n538) );
  NAND2_X1 U589 ( .A1(G113), .A2(n891), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G101), .A2(n895), .ZN(n534) );
  XNOR2_X1 U592 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X2 U594 ( .A(KEYINPUT64), .B(n539), .ZN(G160) );
  INV_X1 U595 ( .A(G651), .ZN(n544) );
  NOR2_X1 U596 ( .A1(G543), .A2(n544), .ZN(n541) );
  XNOR2_X1 U597 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n541), .B(n540), .ZN(n656) );
  NAND2_X1 U599 ( .A1(G64), .A2(n656), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  NAND2_X1 U601 ( .A1(G52), .A2(n657), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G77), .A2(n652), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G90), .A2(n653), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT66), .B(n550), .Z(G301) );
  INV_X1 U609 ( .A(G301), .ZN(G171) );
  NAND2_X1 U610 ( .A1(G72), .A2(n652), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G85), .A2(n653), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G60), .A2(n656), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G47), .A2(n657), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U616 ( .A1(n556), .A2(n555), .ZN(G290) );
  XNOR2_X1 U617 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U618 ( .A(G2451), .B(G2454), .Z(n558) );
  XNOR2_X1 U619 ( .A(G2430), .B(KEYINPUT108), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(n559), .B(G2446), .Z(n561) );
  XNOR2_X1 U622 ( .A(G1341), .B(G1348), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n561), .B(n560), .ZN(n565) );
  XOR2_X1 U624 ( .A(G2438), .B(G2427), .Z(n563) );
  XNOR2_X1 U625 ( .A(G2443), .B(G2435), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U627 ( .A(n565), .B(n564), .Z(n566) );
  AND2_X1 U628 ( .A1(G14), .A2(n566), .ZN(G401) );
  AND2_X1 U629 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  NAND2_X1 U632 ( .A1(G63), .A2(n656), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G51), .A2(n657), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT6), .B(n569), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G89), .A2(n653), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT74), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G76), .A2(n652), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT5), .B(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT75), .B(n575), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT7), .B(n578), .Z(G168) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G65), .A2(n656), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G53), .A2(n657), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT68), .B(n581), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G78), .A2(n652), .ZN(n582) );
  XNOR2_X1 U651 ( .A(KEYINPUT67), .B(n582), .ZN(n583) );
  NOR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n653), .A2(G91), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(G299) );
  XOR2_X1 U655 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n589) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n587) );
  XOR2_X1 U657 ( .A(n587), .B(KEYINPUT10), .Z(n925) );
  NAND2_X1 U658 ( .A1(G567), .A2(n925), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n589), .B(n588), .ZN(G234) );
  NAND2_X1 U660 ( .A1(n653), .A2(G81), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT12), .B(n590), .Z(n593) );
  NAND2_X1 U662 ( .A1(n652), .A2(G68), .ZN(n591) );
  XOR2_X1 U663 ( .A(n591), .B(KEYINPUT72), .Z(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G56), .A2(n656), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n597), .B(KEYINPUT14), .ZN(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT71), .B(n598), .ZN(n599) );
  NOR2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n657), .A2(G43), .ZN(n601) );
  INV_X1 U670 ( .A(G860), .ZN(n614) );
  OR2_X1 U671 ( .A1(n1006), .A2(n614), .ZN(G153) );
  NAND2_X1 U672 ( .A1(G301), .A2(G868), .ZN(n611) );
  NAND2_X1 U673 ( .A1(G66), .A2(n656), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G54), .A2(n657), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G79), .A2(n652), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G92), .A2(n653), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U680 ( .A(n609), .B(KEYINPUT15), .Z(n1012) );
  INV_X1 U681 ( .A(n1012), .ZN(n849) );
  INV_X1 U682 ( .A(G868), .ZN(n673) );
  NAND2_X1 U683 ( .A1(n849), .A2(n673), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G284) );
  NOR2_X1 U685 ( .A1(G286), .A2(n673), .ZN(n613) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U688 ( .A1(G559), .A2(n614), .ZN(n615) );
  XNOR2_X1 U689 ( .A(KEYINPUT76), .B(n615), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n616), .A2(n1012), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT16), .B(n617), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G868), .A2(n1006), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G868), .A2(n1012), .ZN(n618) );
  NOR2_X1 U694 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U695 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G111), .A2(n891), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G99), .A2(n895), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT77), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G135), .A2(n518), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n517), .A2(G123), .ZN(n626) );
  XOR2_X1 U703 ( .A(KEYINPUT18), .B(n626), .Z(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U705 ( .A(KEYINPUT78), .B(n629), .Z(n951) );
  XOR2_X1 U706 ( .A(n951), .B(G2096), .Z(n631) );
  XNOR2_X1 U707 ( .A(G2100), .B(KEYINPUT79), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U709 ( .A1(G49), .A2(n657), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U712 ( .A(KEYINPUT83), .B(n634), .Z(n635) );
  NOR2_X1 U713 ( .A1(n656), .A2(n635), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n636), .A2(G87), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G75), .A2(n652), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G88), .A2(n653), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G62), .A2(n656), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G50), .A2(n657), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(G166) );
  INV_X1 U723 ( .A(G166), .ZN(G303) );
  NAND2_X1 U724 ( .A1(G86), .A2(n653), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G61), .A2(n656), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G73), .A2(n652), .ZN(n647) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n647), .Z(n648) );
  NOR2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n657), .A2(G48), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G80), .A2(n652), .ZN(n655) );
  NAND2_X1 U733 ( .A1(G93), .A2(n653), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n662) );
  NAND2_X1 U735 ( .A1(G67), .A2(n656), .ZN(n659) );
  NAND2_X1 U736 ( .A1(G55), .A2(n657), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT81), .B(n660), .Z(n661) );
  NOR2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT82), .B(n663), .Z(n845) );
  XOR2_X1 U741 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n664) );
  XNOR2_X1 U742 ( .A(G288), .B(n664), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n845), .B(n665), .ZN(n667) );
  XOR2_X1 U744 ( .A(G299), .B(G303), .Z(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n668), .B(G305), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(G290), .ZN(n848) );
  XNOR2_X1 U748 ( .A(n1006), .B(KEYINPUT80), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n1012), .A2(G559), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n671), .B(n670), .ZN(n843) );
  XOR2_X1 U751 ( .A(n848), .B(n843), .Z(n672) );
  NOR2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n675) );
  NOR2_X1 U753 ( .A1(n845), .A2(G868), .ZN(n674) );
  NOR2_X1 U754 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NAND2_X1 U761 ( .A1(G120), .A2(G108), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G69), .A2(n681), .ZN(n846) );
  NAND2_X1 U764 ( .A1(G567), .A2(n846), .ZN(n682) );
  XNOR2_X1 U765 ( .A(n682), .B(KEYINPUT85), .ZN(n687) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n683) );
  XNOR2_X1 U767 ( .A(KEYINPUT22), .B(n683), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n684), .A2(G96), .ZN(n685) );
  OR2_X1 U769 ( .A1(G218), .A2(n685), .ZN(n847) );
  AND2_X1 U770 ( .A1(G2106), .A2(n847), .ZN(n686) );
  NOR2_X1 U771 ( .A1(n687), .A2(n686), .ZN(G319) );
  INV_X1 U772 ( .A(G319), .ZN(n917) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n917), .A2(n688), .ZN(n842) );
  NAND2_X1 U775 ( .A1(n842), .A2(G36), .ZN(G176) );
  NOR2_X1 U776 ( .A1(n710), .A2(n711), .ZN(n834) );
  NAND2_X1 U777 ( .A1(n895), .A2(G105), .ZN(n690) );
  XNOR2_X1 U778 ( .A(KEYINPUT90), .B(KEYINPUT38), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n690), .B(n689), .ZN(n697) );
  NAND2_X1 U780 ( .A1(G117), .A2(n891), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G141), .A2(n518), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U783 ( .A1(G129), .A2(n517), .ZN(n693) );
  XNOR2_X1 U784 ( .A(KEYINPUT89), .B(n693), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U787 ( .A(KEYINPUT91), .B(n698), .Z(n903) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n903), .ZN(n707) );
  NAND2_X1 U789 ( .A1(G107), .A2(n891), .ZN(n700) );
  NAND2_X1 U790 ( .A1(G131), .A2(n518), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n895), .A2(G95), .ZN(n701) );
  XOR2_X1 U793 ( .A(KEYINPUT88), .B(n701), .Z(n702) );
  NOR2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n517), .A2(G119), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n905) );
  NAND2_X1 U797 ( .A1(G1991), .A2(n905), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n949) );
  NAND2_X1 U799 ( .A1(n834), .A2(n949), .ZN(n708) );
  XOR2_X1 U800 ( .A(KEYINPUT92), .B(n708), .Z(n825) );
  XOR2_X1 U801 ( .A(n825), .B(KEYINPUT93), .Z(n808) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n709) );
  XNOR2_X1 U803 ( .A(KEYINPUT24), .B(n709), .ZN(n716) );
  INV_X1 U804 ( .A(n710), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n764), .A2(G8), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n714), .B(n713), .ZN(n715) );
  INV_X1 U807 ( .A(n799), .ZN(n785) );
  NAND2_X1 U808 ( .A1(n716), .A2(n785), .ZN(n784) );
  INV_X1 U809 ( .A(KEYINPUT27), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n743), .A2(G2072), .ZN(n717) );
  XNOR2_X1 U811 ( .A(n718), .B(n717), .ZN(n738) );
  NAND2_X1 U812 ( .A1(G1956), .A2(n764), .ZN(n737) );
  INV_X1 U813 ( .A(G299), .ZN(n719) );
  AND2_X1 U814 ( .A1(n737), .A2(n719), .ZN(n720) );
  AND2_X1 U815 ( .A1(n738), .A2(n720), .ZN(n721) );
  XNOR2_X1 U816 ( .A(n721), .B(KEYINPUT98), .ZN(n735) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n764), .ZN(n723) );
  NAND2_X1 U818 ( .A1(G2067), .A2(n743), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n849), .A2(n731), .ZN(n730) );
  AND2_X1 U821 ( .A1(n743), .A2(G1996), .ZN(n725) );
  XNOR2_X1 U822 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n764), .A2(G1341), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U825 ( .A1(n1006), .A2(n728), .ZN(n729) );
  NOR2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n733) );
  AND2_X1 U827 ( .A1(n849), .A2(n731), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U830 ( .A(n736), .B(KEYINPUT99), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U832 ( .A1(G299), .A2(n739), .ZN(n740) );
  XNOR2_X1 U833 ( .A(n521), .B(KEYINPUT29), .ZN(n748) );
  XOR2_X1 U834 ( .A(KEYINPUT25), .B(G2078), .Z(n926) );
  NOR2_X1 U835 ( .A1(n926), .A2(n764), .ZN(n742) );
  XNOR2_X1 U836 ( .A(n742), .B(KEYINPUT96), .ZN(n745) );
  NOR2_X1 U837 ( .A1(n743), .A2(G1961), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U839 ( .A(KEYINPUT97), .B(n746), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n755), .A2(G171), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n761) );
  NOR2_X1 U842 ( .A1(n799), .A2(G1966), .ZN(n775) );
  NOR2_X1 U843 ( .A1(n764), .A2(G2084), .ZN(n749) );
  XOR2_X1 U844 ( .A(n749), .B(KEYINPUT95), .Z(n774) );
  INV_X1 U845 ( .A(n774), .ZN(n750) );
  NAND2_X1 U846 ( .A1(G8), .A2(n750), .ZN(n751) );
  NOR2_X1 U847 ( .A1(n775), .A2(n751), .ZN(n753) );
  XNOR2_X1 U848 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U849 ( .A1(G168), .A2(n754), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n755), .A2(G171), .ZN(n756) );
  NOR2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U852 ( .A(KEYINPUT31), .B(n758), .ZN(n759) );
  INV_X1 U853 ( .A(n759), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U855 ( .A(n762), .B(KEYINPUT100), .ZN(n777) );
  AND2_X1 U856 ( .A1(G286), .A2(G8), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n777), .A2(n763), .ZN(n772) );
  INV_X1 U858 ( .A(G8), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n799), .A2(G1971), .ZN(n766) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n764), .ZN(n765) );
  NOR2_X1 U861 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U862 ( .A1(n767), .A2(G303), .ZN(n768) );
  XNOR2_X1 U863 ( .A(n768), .B(KEYINPUT102), .ZN(n769) );
  OR2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U866 ( .A(n773), .B(KEYINPUT32), .ZN(n789) );
  AND2_X1 U867 ( .A1(G8), .A2(n774), .ZN(n776) );
  XNOR2_X1 U868 ( .A(n778), .B(KEYINPUT101), .ZN(n787) );
  NAND2_X1 U869 ( .A1(n789), .A2(n787), .ZN(n781) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n782), .A2(n799), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n806) );
  XNOR2_X1 U875 ( .A(G1981), .B(G305), .ZN(n998) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  NAND2_X1 U877 ( .A1(n1004), .A2(n785), .ZN(n791) );
  INV_X1 U878 ( .A(n791), .ZN(n786) );
  AND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n788) );
  AND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n795) );
  NOR2_X1 U881 ( .A1(G1976), .A2(G288), .ZN(n796) );
  NOR2_X1 U882 ( .A1(G1971), .A2(G303), .ZN(n790) );
  NOR2_X1 U883 ( .A1(n796), .A2(n790), .ZN(n1015) );
  OR2_X1 U884 ( .A1(n791), .A2(n1015), .ZN(n793) );
  INV_X1 U885 ( .A(KEYINPUT33), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n802) );
  NAND2_X1 U888 ( .A1(KEYINPUT33), .A2(n796), .ZN(n797) );
  XOR2_X1 U889 ( .A(KEYINPUT103), .B(n797), .Z(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n800), .B(KEYINPUT104), .ZN(n801) );
  NOR2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U893 ( .A(n803), .B(KEYINPUT105), .ZN(n804) );
  NOR2_X1 U894 ( .A1(n998), .A2(n804), .ZN(n805) );
  NOR2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n821) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n1003) );
  NAND2_X1 U898 ( .A1(n1003), .A2(n834), .ZN(n809) );
  XOR2_X1 U899 ( .A(KEYINPUT87), .B(n809), .Z(n819) );
  XOR2_X1 U900 ( .A(G2067), .B(KEYINPUT37), .Z(n832) );
  NAND2_X1 U901 ( .A1(G104), .A2(n895), .ZN(n811) );
  NAND2_X1 U902 ( .A1(G140), .A2(n518), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U904 ( .A(KEYINPUT34), .B(n812), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G116), .A2(n891), .ZN(n814) );
  NAND2_X1 U906 ( .A1(G128), .A2(n517), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT35), .B(n815), .Z(n816) );
  NOR2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U910 ( .A(KEYINPUT36), .B(n818), .Z(n914) );
  AND2_X1 U911 ( .A1(n832), .A2(n914), .ZN(n950) );
  NAND2_X1 U912 ( .A1(n950), .A2(n834), .ZN(n822) );
  AND2_X1 U913 ( .A1(n819), .A2(n822), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n838) );
  INV_X1 U915 ( .A(n822), .ZN(n831) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n905), .ZN(n954) );
  NOR2_X1 U918 ( .A1(n823), .A2(n954), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n827) );
  NOR2_X1 U920 ( .A1(n903), .A2(G1996), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n826), .B(KEYINPUT106), .ZN(n947) );
  NOR2_X1 U922 ( .A1(n827), .A2(n947), .ZN(n828) );
  XNOR2_X1 U923 ( .A(KEYINPUT39), .B(n828), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n834), .A2(n829), .ZN(n830) );
  OR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n836) );
  NOR2_X1 U926 ( .A1(n832), .A2(n914), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(n833), .Z(n968) );
  NAND2_X1 U928 ( .A1(n968), .A2(n834), .ZN(n835) );
  AND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U931 ( .A(n839), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n925), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G188) );
  XNOR2_X1 U937 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  NOR2_X1 U939 ( .A1(n843), .A2(G860), .ZN(n844) );
  XOR2_X1 U940 ( .A(n845), .B(n844), .Z(G145) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  XOR2_X1 U945 ( .A(KEYINPUT114), .B(n848), .Z(n851) );
  XOR2_X1 U946 ( .A(n849), .B(G286), .Z(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U948 ( .A(n1006), .B(G171), .Z(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  NOR2_X1 U950 ( .A1(G37), .A2(n854), .ZN(G397) );
  XOR2_X1 U951 ( .A(G2100), .B(G2096), .Z(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(G2678), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2090), .Z(n858) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U960 ( .A(G1976), .B(G1961), .Z(n864) );
  XNOR2_X1 U961 ( .A(G1981), .B(G1966), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n869) );
  XOR2_X1 U963 ( .A(G1991), .B(G1986), .Z(n867) );
  INV_X1 U964 ( .A(G1996), .ZN(n865) );
  XOR2_X1 U965 ( .A(n865), .B(G1971), .Z(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U968 ( .A(KEYINPUT109), .B(G2474), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n873) );
  XOR2_X1 U970 ( .A(G1956), .B(KEYINPUT41), .Z(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U972 ( .A1(G124), .A2(n517), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n874), .B(KEYINPUT110), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G100), .A2(n895), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G112), .A2(n891), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G136), .A2(n518), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT111), .B(n882), .Z(G162) );
  NAND2_X1 U982 ( .A1(G103), .A2(n895), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G139), .A2(n518), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n891), .A2(G115), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n885), .B(KEYINPUT112), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G127), .A2(n517), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n958) );
  NAND2_X1 U991 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G130), .A2(n517), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U994 ( .A1(G106), .A2(n895), .ZN(n898) );
  NAND2_X1 U995 ( .A1(G142), .A2(n518), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT45), .B(n899), .Z(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n958), .B(n902), .ZN(n913) );
  XNOR2_X1 U1000 ( .A(G162), .B(G160), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n905), .B(KEYINPUT46), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G164), .B(n951), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n917), .ZN(n922) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1013 ( .A(KEYINPUT115), .B(n918), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n919), .B(KEYINPUT49), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G397), .A2(n920), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1017 ( .A1(n923), .A2(G395), .ZN(n924) );
  XOR2_X1 U1018 ( .A(n924), .B(KEYINPUT116), .Z(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  INV_X1 U1021 ( .A(n925), .ZN(G223) );
  XOR2_X1 U1022 ( .A(G32), .B(G1996), .Z(n938) );
  XOR2_X1 U1023 ( .A(n926), .B(G27), .Z(n932) );
  XOR2_X1 U1024 ( .A(G2067), .B(G26), .Z(n927) );
  XNOR2_X1 U1025 ( .A(KEYINPUT121), .B(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT122), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n936) );
  XOR2_X1 U1030 ( .A(G1991), .B(G25), .Z(n933) );
  NAND2_X1 U1031 ( .A1(n933), .A2(G28), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(KEYINPUT120), .B(n934), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n939), .B(KEYINPUT53), .ZN(n942) );
  XOR2_X1 U1036 ( .A(G2084), .B(KEYINPUT54), .Z(n940) );
  XNOR2_X1 U1037 ( .A(G34), .B(n940), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G35), .B(G2090), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n1028) );
  NAND2_X1 U1041 ( .A1(KEYINPUT55), .A2(n1028), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n945), .ZN(n1027) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1045 ( .A(KEYINPUT51), .B(n948), .Z(n966) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(G2084), .B(G160), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT118), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n964) );
  XOR2_X1 U1052 ( .A(n958), .B(KEYINPUT119), .Z(n959) );
  XOR2_X1 U1053 ( .A(G2072), .B(n959), .Z(n961) );
  XOR2_X1 U1054 ( .A(G164), .B(G2078), .Z(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT50), .B(n962), .Z(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT52), .B(n969), .ZN(n971) );
  INV_X1 U1061 ( .A(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n973), .B(G4), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G1956), .B(G20), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(KEYINPUT124), .B(G1341), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G19), .B(n978), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT60), .B(n981), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G21), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G1961), .B(G5), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(G23), .B(G1976), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G1986), .B(KEYINPUT125), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n988), .B(G24), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(n994), .B(KEYINPUT126), .Z(n995) );
  XNOR2_X1 U1087 ( .A(KEYINPUT61), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n996), .ZN(n1022) );
  XOR2_X1 U1089 ( .A(G16), .B(KEYINPUT56), .Z(n1020) );
  XOR2_X1 U1090 ( .A(G168), .B(G1966), .Z(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1092 ( .A(KEYINPUT57), .B(n999), .Z(n1011) );
  XOR2_X1 U1093 ( .A(G1956), .B(G299), .Z(n1001) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n1000) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(G1341), .B(n1006), .Z(n1007) );
  XNOR2_X1 U1099 ( .A(KEYINPUT123), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(n1012), .B(G1348), .Z(n1014) );
  XOR2_X1 U1103 ( .A(G171), .B(G1961), .Z(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT127), .B(n1023), .Z(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1032) );
  INV_X1 U1112 ( .A(n1028), .ZN(n1030) );
  NOR2_X1 U1113 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
endmodule

