//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT2), .A3(G113), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n189), .A2(new_n191), .B1(new_n187), .B2(new_n188), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(KEYINPUT68), .A3(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT69), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT69), .B1(new_n192), .B2(new_n199), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT0), .A3(G128), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT0), .B(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT11), .A2(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT64), .A2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n212), .A2(new_n213), .A3(new_n217), .A4(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT11), .A2(G134), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n213), .B1(new_n220), .B2(new_n211), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AOI211_X1 g037(.A(G131), .B(new_n221), .C1(new_n216), .C2(new_n218), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n208), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n219), .A2(new_n209), .A3(new_n222), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT64), .A2(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT64), .A2(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(G131), .C1(new_n230), .C2(new_n211), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(G128), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n234), .B(new_n236), .C1(KEYINPUT1), .C2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(new_n232), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n225), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n225), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT66), .B(new_n208), .C1(new_n223), .C2(new_n224), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n203), .B(new_n244), .C1(new_n249), .C2(KEYINPUT30), .ZN(new_n250));
  INV_X1    g064(.A(new_n203), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n225), .A2(new_n251), .A3(new_n243), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT31), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n250), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n252), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n252), .B1(new_n249), .B2(new_n251), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n260), .B(new_n262), .C1(new_n257), .C2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(G472), .A2(G902), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n270), .A2(KEYINPUT32), .A3(new_n271), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n225), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n203), .B1(new_n279), .B2(new_n245), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n263), .B1(new_n280), .B2(new_n252), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n264), .A2(KEYINPUT29), .A3(new_n257), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n217), .B1(new_n229), .B2(new_n213), .ZN(new_n286));
  INV_X1    g100(.A(new_n218), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n222), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n226), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT66), .B1(new_n290), .B2(new_n208), .ZN(new_n291));
  INV_X1    g105(.A(new_n248), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n243), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n203), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n267), .B1(new_n294), .B2(new_n252), .ZN(new_n295));
  INV_X1    g109(.A(new_n257), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n265), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n285), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n257), .B1(new_n250), .B2(new_n252), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n284), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n277), .B1(new_n301), .B2(G472), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n266), .A2(new_n268), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n303), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n250), .A2(new_n252), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n296), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n283), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G472), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(KEYINPUT72), .A3(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n275), .B(new_n276), .C1(new_n302), .C2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT24), .B(G110), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n240), .A2(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n196), .A2(G128), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n317));
  INV_X1    g131(.A(new_n313), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n314), .C1(new_n318), .C2(KEYINPUT23), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT75), .B(G110), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n321), .B2(KEYINPUT76), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(KEYINPUT76), .B2(new_n321), .ZN(new_n323));
  AND2_X1   g137(.A1(KEYINPUT74), .A2(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(KEYINPUT74), .A2(G125), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G140), .B1(new_n324), .B2(new_n325), .ZN(new_n331));
  OR2_X1    g145(.A1(G125), .A2(G140), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n330), .B(G146), .C1(new_n333), .C2(new_n328), .ZN(new_n334));
  XNOR2_X1  g148(.A(G125), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n233), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n323), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n233), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n319), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n343), .B2(new_n319), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n312), .A2(new_n315), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n341), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n337), .A2(new_n347), .A3(new_n352), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n356), .B2(KEYINPUT77), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n359), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n354), .A2(new_n361), .A3(new_n355), .A4(new_n357), .ZN(new_n362));
  INV_X1    g176(.A(G217), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(G234), .B2(new_n278), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n354), .A2(new_n355), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n207), .A2(new_n327), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n239), .A2(new_n241), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n326), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n350), .A2(G224), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n374), .B(KEYINPUT85), .Z(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n192), .A2(new_n199), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(G107), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT79), .B(G101), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(G104), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n387), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n388), .A2(new_n390), .B1(G101), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n188), .B1(new_n194), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n197), .A2(new_n198), .ZN(new_n396));
  INV_X1    g210(.A(new_n194), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n395), .B1(new_n398), .B2(new_n394), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT82), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(new_n395), .C1(new_n398), .C2(new_n394), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n381), .A2(new_n393), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT4), .A3(G101), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n388), .B2(new_n390), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(G101), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n203), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n403), .A2(new_n410), .A3(new_n412), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n403), .B2(new_n410), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n417), .A2(KEYINPUT84), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT84), .B1(new_n417), .B2(new_n419), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n376), .B(new_n416), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n374), .A2(KEYINPUT7), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n370), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n373), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n370), .B(new_n372), .C1(new_n424), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n392), .A2(G101), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n404), .B2(new_n389), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n381), .A2(new_n430), .A3(new_n400), .A4(new_n402), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n412), .B(KEYINPUT8), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n381), .A2(new_n399), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n393), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n428), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n415), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n422), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT87), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n422), .A2(new_n436), .ZN(new_n440));
  INV_X1    g254(.A(new_n437), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n422), .A2(new_n443), .A3(new_n436), .A4(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G478), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT15), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT96), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n193), .A3(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT95), .ZN(new_n453));
  INV_X1    g267(.A(G122), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n454), .B2(G116), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n455), .C1(new_n193), .C2(G122), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n452), .A2(KEYINPUT95), .ZN(new_n457));
  OAI21_X1  g271(.A(G107), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G116), .B(G122), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n385), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n235), .A2(G128), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n240), .A2(G143), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT94), .ZN(new_n466));
  AOI21_X1  g280(.A(G134), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n465), .A2(G134), .A3(new_n466), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n458), .B(new_n460), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT9), .B(G234), .Z(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT78), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(G217), .A3(new_n350), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n467), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n459), .B(new_n385), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n462), .B1(new_n461), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n461), .A2(new_n476), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT93), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n461), .A2(new_n480), .A3(new_n476), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n474), .B(new_n475), .C1(new_n230), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n473), .B1(new_n469), .B2(new_n483), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n278), .B(new_n450), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT97), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n278), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n449), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G234), .A2(G237), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n493), .A2(G952), .A3(new_n350), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n493), .A2(G902), .A3(G953), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT21), .B(G898), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n430), .A2(new_n371), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT80), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n393), .A2(new_n242), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT80), .B1(new_n430), .B2(new_n371), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT81), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n430), .A2(new_n371), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n290), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT12), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n430), .A2(new_n371), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n409), .A2(new_n208), .B1(new_n509), .B2(KEYINPUT10), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n223), .A2(new_n224), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n502), .A2(new_n512), .A3(new_n503), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G110), .B(G140), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n350), .A2(G227), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n506), .A2(new_n519), .A3(new_n290), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n508), .A2(new_n514), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n511), .B1(new_n510), .B2(new_n513), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G469), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n278), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n508), .A2(new_n514), .A3(new_n520), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n522), .A2(new_n523), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n518), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n533), .A3(G469), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G221), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n471), .B2(new_n278), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n253), .A2(G214), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n235), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n209), .A3(new_n540), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n540), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT17), .A3(G131), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n334), .A2(new_n340), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n382), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT89), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(KEYINPUT18), .A3(G131), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n331), .A2(new_n332), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n336), .B1(new_n556), .B2(new_n233), .ZN(new_n557));
  NAND2_X1  g371(.A1(KEYINPUT18), .A2(G131), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n545), .A2(new_n540), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n551), .A2(new_n554), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n543), .A2(new_n546), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n335), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n233), .B(new_n564), .C1(new_n556), .C2(new_n563), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n334), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n553), .B1(new_n566), .B2(new_n560), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n539), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT91), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n560), .ZN(new_n571));
  INV_X1    g385(.A(new_n553), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n551), .A2(new_n554), .A3(new_n560), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT90), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n576), .A2(new_n577), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G475), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n551), .A2(new_n560), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n553), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n551), .A2(KEYINPUT92), .A3(new_n560), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n574), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n582), .B1(new_n588), .B2(new_n278), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n581), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n498), .A2(new_n535), .A3(new_n538), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n447), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n310), .A2(new_n369), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n389), .ZN(G3));
  NOR2_X1   g408(.A1(new_n269), .A2(new_n257), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n261), .B1(new_n250), .B2(new_n258), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n250), .A2(new_n261), .A3(new_n258), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n598), .B2(G902), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(KEYINPUT98), .B1(new_n271), .B2(new_n270), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n601), .B(G472), .C1(new_n598), .C2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n535), .A2(new_n538), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n368), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n606));
  INV_X1    g420(.A(new_n446), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n606), .B(new_n438), .C1(new_n442), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n438), .A2(new_n606), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n437), .B1(new_n422), .B2(new_n436), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n576), .A2(new_n577), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n578), .A2(new_n580), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n561), .B1(new_n585), .B2(new_n586), .ZN(new_n616));
  OAI21_X1  g430(.A(G475), .B1(new_n616), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n497), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n469), .A2(new_n483), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n622), .B2(KEYINPUT100), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n485), .B2(new_n486), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n622), .B(new_n484), .C1(KEYINPUT100), .C2(new_n620), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(G478), .A3(new_n625), .ZN(new_n626));
  MUX2_X1   g440(.A(new_n278), .B(new_n490), .S(new_n448), .Z(new_n627));
  AND2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n619), .A3(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n605), .A2(new_n612), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n634), .B(G475), .C1(new_n616), .C2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n576), .B(new_n577), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n492), .A2(new_n636), .A3(new_n637), .A4(new_n619), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n638), .A2(new_n608), .A3(new_n611), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n605), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR2_X1   g458(.A1(new_n597), .A2(new_n596), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n296), .B1(new_n295), .B2(new_n265), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT98), .B1(new_n647), .B2(new_n308), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n602), .A3(new_n272), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n491), .A2(new_n487), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(KEYINPUT97), .B2(new_n487), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n590), .A2(new_n651), .A3(new_n619), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n603), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n348), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n366), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n365), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n653), .A2(new_n446), .A3(new_n445), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n649), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT103), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT37), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(new_n612), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n494), .B1(new_n495), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n492), .A2(new_n636), .A3(new_n637), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n657), .A2(new_n535), .A3(new_n538), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n310), .A2(new_n663), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  XOR2_X1   g485(.A(new_n665), .B(KEYINPUT39), .Z(new_n672));
  NAND3_X1  g486(.A1(new_n535), .A2(new_n538), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n445), .B(KEYINPUT38), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n296), .B1(new_n250), .B2(new_n252), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n280), .A2(new_n252), .A3(new_n296), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n278), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n275), .A2(new_n276), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n618), .A2(new_n492), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n607), .A3(new_n657), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n674), .A2(new_n675), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NAND3_X1  g498(.A1(new_n628), .A2(new_n618), .A3(new_n666), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n310), .A2(new_n663), .A3(new_n669), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NOR2_X1   g502(.A1(new_n612), .A2(new_n629), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n521), .A2(new_n524), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n526), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n691), .A2(G902), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n525), .A2(new_n692), .A3(new_n526), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n538), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n310), .A2(new_n689), .A3(new_n369), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT105), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n699), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n310), .A2(new_n369), .A3(new_n639), .A4(new_n698), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NOR2_X1   g518(.A1(new_n612), .A2(new_n697), .ZN(new_n705));
  INV_X1    g519(.A(new_n657), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n652), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n310), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NOR2_X1   g523(.A1(new_n612), .A2(new_n681), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n308), .B1(new_n270), .B2(new_n278), .ZN(new_n711));
  INV_X1    g525(.A(new_n271), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n296), .B1(new_n281), .B2(new_n265), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n645), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n711), .A2(new_n368), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n710), .A2(new_n619), .A3(new_n715), .A4(new_n698), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NOR3_X1   g531(.A1(new_n711), .A2(new_n706), .A3(new_n714), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n705), .A2(new_n686), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT32), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n721), .B(new_n712), .C1(new_n645), .C2(new_n646), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT108), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n301), .A2(new_n277), .A3(G472), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT72), .B1(new_n307), .B2(new_n308), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n272), .A2(new_n721), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n531), .B2(new_n533), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT106), .B1(new_n530), .B2(new_n517), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n526), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n527), .A2(new_n529), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n538), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n439), .A2(new_n442), .A3(new_n446), .A4(new_n444), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n685), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n369), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n310), .A2(new_n369), .A3(new_n686), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n739), .A2(KEYINPUT107), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NAND4_X1  g558(.A1(new_n310), .A2(new_n369), .A3(new_n667), .A4(new_n738), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NAND2_X1  g560(.A1(new_n628), .A2(new_n590), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n649), .A2(new_n657), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT44), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n730), .A2(new_n731), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT45), .B1(new_n531), .B2(new_n533), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n526), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n528), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n527), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n538), .B(new_n672), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n735), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n751), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  INV_X1    g576(.A(new_n310), .ZN(new_n763));
  INV_X1    g577(.A(new_n735), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n368), .A3(new_n686), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n538), .B1(new_n757), .B2(new_n758), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT47), .B(new_n538), .C1(new_n757), .C2(new_n758), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT109), .B(G140), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G42));
  INV_X1    g586(.A(new_n680), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n697), .A2(new_n735), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n369), .A3(new_n494), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n775), .A2(new_n618), .A3(new_n628), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT114), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n749), .A2(new_n494), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n774), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n777), .B1(new_n718), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n780), .A2(new_n715), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n675), .A2(new_n446), .A3(new_n697), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(KEYINPUT50), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n780), .A2(new_n715), .A3(new_n764), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g605(.A(new_n696), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n768), .B(new_n769), .C1(new_n538), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n782), .A2(new_n789), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n782), .A2(new_n789), .A3(KEYINPUT51), .A4(new_n795), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n781), .A2(new_n369), .A3(new_n728), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT48), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n783), .A2(new_n705), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n626), .B(new_n627), .C1(new_n581), .C2(new_n589), .ZN(new_n805));
  OAI211_X1 g619(.A(G952), .B(new_n350), .C1(new_n775), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n798), .A2(new_n799), .A3(new_n801), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n636), .A2(new_n651), .A3(new_n637), .A4(new_n666), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n668), .A2(new_n735), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n310), .A2(new_n810), .B1(new_n736), .B2(new_n718), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n745), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT110), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n745), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n600), .A2(new_n592), .A3(new_n602), .A4(new_n657), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n492), .A2(new_n615), .A3(new_n617), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n497), .B1(new_n818), .B2(new_n805), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n819), .A2(new_n446), .A3(new_n445), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n600), .A2(new_n820), .A3(new_n602), .A4(new_n604), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n699), .A2(new_n703), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n593), .A2(new_n708), .A3(new_n716), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n743), .A2(new_n816), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n734), .A2(new_n657), .A3(new_n665), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n710), .A2(new_n680), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n670), .A2(new_n687), .A3(new_n719), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT52), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n670), .A2(new_n719), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n687), .A4(new_n827), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n835), .B2(KEYINPUT111), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n830), .B(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n825), .B2(new_n829), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n811), .A2(new_n745), .A3(new_n814), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n814), .B1(new_n811), .B2(new_n745), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n593), .A2(new_n708), .A3(new_n716), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n703), .A2(new_n821), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n273), .B1(new_n270), .B2(new_n271), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n722), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n368), .B(new_n697), .C1(new_n847), .C2(new_n726), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n659), .B1(new_n848), .B2(new_n689), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n743), .A4(new_n835), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n840), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n838), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n808), .A2(new_n839), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n792), .A2(KEYINPUT49), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n369), .A2(new_n446), .A3(new_n538), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n859), .A2(new_n747), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n773), .C1(KEYINPUT49), .C2(new_n792), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n857), .A2(new_n858), .B1(new_n675), .B2(new_n862), .ZN(G75));
  NOR2_X1   g677(.A1(new_n854), .A2(new_n278), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(G210), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n376), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  XOR2_X1   g682(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n869));
  AND3_X1   g683(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n350), .A2(G952), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(G51));
  AND3_X1   g688(.A1(new_n864), .A2(new_n753), .A3(new_n755), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n840), .A2(new_n853), .A3(KEYINPUT54), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n855), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n528), .B(KEYINPUT117), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT57), .Z(new_n879));
  AOI21_X1  g693(.A(new_n691), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n879), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n855), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT118), .B1(new_n884), .B2(new_n691), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n873), .B1(new_n882), .B2(new_n885), .ZN(G54));
  NAND3_X1  g700(.A1(new_n864), .A2(KEYINPUT58), .A3(G475), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n568), .A2(new_n575), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n873), .ZN(G60));
  NAND2_X1  g705(.A1(new_n624), .A2(new_n625), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT119), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n448), .A2(new_n278), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n894), .B(new_n895), .Z(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n877), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n873), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n896), .B1(new_n839), .B2(new_n856), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n893), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n840), .A2(new_n853), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n354), .A2(new_n355), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n873), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n840), .A2(new_n853), .A3(new_n655), .A4(new_n906), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT61), .B1(new_n909), .B2(KEYINPUT122), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(G66));
  INV_X1    g729(.A(G224), .ZN(new_n916));
  OAI21_X1  g730(.A(G953), .B1(new_n496), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n824), .B2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n866), .B1(G898), .B2(new_n350), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n918), .B(new_n920), .ZN(G69));
  NAND3_X1  g735(.A1(new_n831), .A2(new_n683), .A3(new_n687), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n770), .B1(new_n760), .B2(new_n751), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n673), .B1(new_n805), .B2(new_n818), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n310), .A2(new_n369), .A3(new_n764), .A4(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n926), .B(new_n928), .C1(KEYINPUT62), .C2(new_n922), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n350), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n244), .B1(new_n249), .B2(KEYINPUT30), .ZN(new_n931));
  INV_X1    g745(.A(new_n564), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n333), .B2(KEYINPUT19), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n930), .A2(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n936), .A2(new_n935), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n728), .A2(new_n369), .A3(new_n710), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n745), .B1(new_n939), .B2(new_n759), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n926), .A2(new_n687), .A3(new_n831), .A4(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n743), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n350), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n664), .A2(G953), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(KEYINPUT125), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n934), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n937), .B(new_n938), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n944), .A2(new_n945), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n947), .A3(new_n946), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n938), .B1(new_n955), .B2(new_n937), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n951), .A2(new_n956), .ZN(G72));
  INV_X1    g771(.A(new_n676), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n925), .A2(new_n929), .A3(new_n850), .ZN(new_n959));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT127), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n942), .A2(new_n943), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n965), .B2(new_n824), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n305), .A2(new_n257), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n900), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n958), .A3(new_n961), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n837), .A2(new_n970), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n964), .A2(new_n969), .A3(new_n971), .ZN(G57));
endmodule


