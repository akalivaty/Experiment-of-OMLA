//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G234));
  NAND2_X1  g025(.A1(new_n447), .A2(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT70), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n467), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n474), .B2(new_n476), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  INV_X1    g058(.A(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n477), .A2(new_n467), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n477), .A2(KEYINPUT72), .A3(new_n478), .A4(new_n467), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n485), .A2(new_n478), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n478), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n491), .A2(G124), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n478), .A3(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n470), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n478), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n477), .A2(new_n467), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n477), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  AND2_X1   g093(.A1(G75), .A2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n511), .B2(new_n513), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI211_X1 g098(.A(G88), .B(new_n517), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI21_X1  g100(.A(G543), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n520), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  OAI211_X1 g103(.A(G51), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n529));
  OAI211_X1 g104(.A(G89), .B(new_n517), .C1(new_n522), .C2(new_n523), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  AND2_X1   g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n531), .A2(new_n535), .A3(G63), .A4(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n529), .A2(new_n530), .A3(new_n536), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n542), .A2(new_n526), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n514), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n531), .A2(new_n535), .A3(G64), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n541), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n545), .A2(new_n541), .A3(new_n549), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n531), .A2(new_n535), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n546), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n559), .A2(new_n526), .B1(new_n543), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n558), .A2(G860), .A3(new_n562), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n533), .A2(new_n534), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT76), .B(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n543), .ZN(new_n577));
  OAI211_X1 g152(.A(G53), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  NOR3_X1   g158(.A1(new_n533), .A2(new_n534), .A3(new_n532), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT74), .B1(new_n515), .B2(new_n516), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(G651), .ZN(new_n588));
  AOI21_X1  g163(.A(G74), .B1(new_n531), .B2(new_n535), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT78), .B1(new_n589), .B2(new_n510), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g166(.A(G49), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n592));
  OAI211_X1 g167(.A(G87), .B(new_n517), .C1(new_n522), .C2(new_n523), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(G288));
  AND2_X1   g170(.A1(new_n517), .A2(G61), .ZN(new_n596));
  AND2_X1   g171(.A1(G73), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n514), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g173(.A(G48), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n599));
  INV_X1    g174(.A(G86), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n543), .ZN(G305));
  INV_X1    g176(.A(new_n526), .ZN(new_n602));
  INV_X1    g177(.A(new_n543), .ZN(new_n603));
  AOI22_X1  g178(.A1(G47), .A2(new_n602), .B1(new_n603), .B2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n555), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n514), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(G290));
  NAND3_X1  g184(.A1(new_n603), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n543), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n602), .A2(G54), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n517), .A2(G66), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT79), .ZN(new_n618));
  OAI21_X1  g193(.A(G651), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n615), .A2(KEYINPUT80), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(KEYINPUT80), .B1(new_n615), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n622), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g198(.A(new_n622), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n581), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(new_n622), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n558), .A2(new_n562), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  MUX2_X1   g207(.A(new_n631), .B(new_n632), .S(G868), .Z(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g210(.A1(new_n480), .A2(new_n467), .A3(new_n469), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2100), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n489), .A2(G135), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n478), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n491), .A2(G123), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT83), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n673), .C1(new_n670), .C2(new_n666), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n666), .A2(new_n668), .A3(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n669), .A2(new_n672), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n674), .B(new_n676), .C1(new_n667), .C2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n682), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n682), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  NOR2_X1   g273(.A1(G5), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G171), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1961), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(G115), .A2(G2104), .ZN(new_n703));
  INV_X1    g278(.A(G127), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n470), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n478), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n706), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G139), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n708), .B(new_n711), .C1(new_n712), .C2(new_n488), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  MUX2_X1   g289(.A(G33), .B(new_n714), .S(G29), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G2072), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n702), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n717), .B1(G2072), .B2(new_n715), .C1(G2090), .C2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G19), .B(new_n631), .S(G16), .Z(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n718), .A2(G27), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G164), .B2(new_n718), .ZN(new_n727));
  INV_X1    g302(.A(G2078), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n482), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n645), .A2(new_n718), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT31), .B(G11), .Z(new_n743));
  INV_X1    g318(.A(G28), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n725), .A2(new_n729), .A3(new_n734), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G2090), .B2(new_n722), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n730), .A2(G20), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT23), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G299), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1956), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n628), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n751), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n718), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n489), .A2(G141), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT26), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n480), .A2(G105), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n764), .B(new_n765), .C1(new_n491), .C2(G129), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(new_n718), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT27), .ZN(new_n769));
  INV_X1    g344(.A(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n489), .A2(G140), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n478), .A2(G116), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n491), .A2(G128), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT88), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n718), .A2(G26), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT28), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  OR4_X1    g358(.A1(new_n723), .A2(new_n760), .A3(new_n771), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G23), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n591), .A2(new_n786), .A3(new_n594), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n591), .B2(new_n594), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n785), .B1(new_n789), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n730), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n730), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G305), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n792), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n790), .A2(new_n791), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n730), .A2(G24), .ZN(new_n806));
  INV_X1    g381(.A(G290), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n730), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1986), .ZN(new_n809));
  OR2_X1    g384(.A1(G25), .A2(G29), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n489), .A2(G131), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT86), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G119), .B2(new_n491), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n718), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n809), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n804), .A2(new_n805), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT36), .Z(new_n823));
  NOR2_X1   g398(.A1(new_n784), .A2(new_n823), .ZN(G311));
  INV_X1    g399(.A(G311), .ZN(G150));
  NAND2_X1  g400(.A1(new_n628), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n556), .A2(G67), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n546), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT93), .B(G93), .Z(new_n832));
  OAI22_X1  g407(.A1(new_n831), .A2(new_n526), .B1(new_n543), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n558), .A3(new_n562), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n557), .A2(new_n546), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n836), .A2(new_n561), .B1(new_n830), .B2(new_n833), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n827), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT94), .B(G860), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n834), .A2(new_n842), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  NAND2_X1  g421(.A1(new_n767), .A2(new_n508), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n762), .A2(new_n766), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G164), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n847), .A2(new_n777), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n777), .B1(new_n847), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n714), .A2(KEYINPUT95), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n714), .A2(KEYINPUT95), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n854), .B(new_n852), .C1(new_n851), .C2(new_n850), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n811), .A2(KEYINPUT97), .A3(new_n815), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT97), .B1(new_n811), .B2(new_n815), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n637), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n489), .A2(G142), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n478), .A2(G118), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT96), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n862), .B2(KEYINPUT96), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n491), .A2(G130), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n816), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n637), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n857), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n860), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n868), .B1(new_n860), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n856), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(new_n853), .A3(new_n855), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n645), .B(new_n482), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n496), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT98), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n883));
  INV_X1    g458(.A(new_n881), .ZN(new_n884));
  AOI211_X1 g459(.A(new_n883), .B(new_n884), .C1(new_n876), .C2(new_n878), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n877), .A2(new_n887), .A3(new_n853), .A4(new_n855), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n873), .B2(new_n874), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n856), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n890), .A3(new_n884), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT100), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT40), .A4(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n882), .B2(new_n885), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n891), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n894), .A2(new_n899), .ZN(G395));
  NAND2_X1  g475(.A1(new_n789), .A2(G305), .ZN(new_n901));
  XNOR2_X1  g476(.A(G290), .B(G303), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n797), .B1(new_n787), .B2(new_n788), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n908), .B2(new_n906), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n622), .B(G299), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n622), .B(new_n581), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n632), .B(new_n838), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n918), .B2(new_n912), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n921));
  OR3_X1    g496(.A1(new_n911), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n919), .B(KEYINPUT102), .C1(new_n918), .C2(new_n912), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n911), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(G868), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n834), .A2(G868), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n926), .B2(new_n930), .ZN(G295));
  AOI21_X1  g506(.A(new_n928), .B1(new_n926), .B2(new_n930), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(new_n906), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n835), .A2(new_n837), .ZN(new_n935));
  OAI21_X1  g510(.A(G168), .B1(new_n551), .B2(new_n552), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n552), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(G286), .A3(new_n550), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n936), .A2(new_n939), .A3(new_n837), .A4(new_n835), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n915), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n838), .B1(new_n936), .B2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n838), .A2(KEYINPUT104), .A3(new_n936), .A4(new_n939), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n914), .A2(new_n916), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n934), .B(new_n943), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n952), .B2(new_n906), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n951), .B1(new_n953), .B2(KEYINPUT105), .ZN(new_n954));
  INV_X1    g529(.A(new_n943), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n947), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n941), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n917), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n893), .B1(new_n958), .B2(new_n934), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n933), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n949), .B1(new_n941), .B2(new_n942), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n956), .A2(new_n915), .A3(new_n941), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n906), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n893), .A3(new_n950), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n954), .A2(new_n961), .A3(new_n933), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT106), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n954), .A2(new_n961), .A3(new_n971), .A4(new_n933), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n968), .B1(new_n974), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n503), .B2(new_n507), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n473), .A2(G40), .A3(new_n479), .A4(new_n481), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n770), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n848), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n777), .A2(G2067), .ZN(new_n984));
  INV_X1    g559(.A(G2067), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n772), .A2(new_n985), .A3(new_n776), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n767), .A2(new_n770), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n981), .B(KEYINPUT108), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n816), .B(new_n818), .Z(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n990), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1986), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n981), .A2(new_n807), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n807), .A2(new_n996), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n981), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT107), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT112), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1006), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n1004), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n976), .C1(new_n503), .C2(new_n507), .ZN(new_n1012));
  INV_X1    g587(.A(new_n980), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n977), .A2(new_n1015), .A3(new_n978), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n977), .B2(new_n978), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1014), .B(new_n1021), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT111), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n976), .C1(new_n503), .C2(new_n507), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(new_n1013), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n977), .A2(new_n1029), .A3(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(G2090), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1003), .B(new_n1011), .C1(new_n1023), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n787), .A2(new_n788), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n977), .B2(new_n980), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G288), .A2(KEYINPUT87), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n591), .A2(new_n786), .A3(new_n594), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G1976), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1037), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1038), .A2(KEYINPUT52), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n603), .A2(G86), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n599), .A4(new_n598), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(new_n1051), .A3(KEYINPUT49), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1043), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1047), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1034), .B1(new_n1045), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1038), .A2(KEYINPUT52), .A3(new_n1044), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1047), .A2(new_n1056), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(KEYINPUT116), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1033), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G286), .A2(G8), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1025), .A2(new_n1028), .A3(new_n740), .A4(new_n1030), .ZN(new_n1067));
  INV_X1    g642(.A(new_n979), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n733), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1003), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1065), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT51), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1066), .A2(new_n1071), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1074), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1065), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1075), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n508), .A2(KEYINPUT114), .A3(new_n1026), .A4(new_n976), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1027), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n980), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G2090), .B1(new_n1088), .B2(KEYINPUT115), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1084), .A2(new_n1087), .A3(new_n1090), .A4(new_n1086), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1023), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G8), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1062), .A2(new_n1081), .A3(new_n1083), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n979), .A2(KEYINPUT109), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n977), .A2(new_n1015), .A3(new_n978), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1021), .B1(new_n1101), .B2(new_n1014), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1022), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n728), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1105), .A2(G2078), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1031), .A2(new_n701), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G301), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G2078), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1111));
  OAI211_X1 g686(.A(G301), .B(new_n1109), .C1(new_n1111), .C2(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1098), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1109), .B1(new_n1111), .B2(KEYINPUT53), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT54), .A3(new_n1112), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT126), .B1(new_n1097), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1023), .A2(new_n1032), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(G8), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT116), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1059), .A2(new_n1060), .A3(KEYINPUT116), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1096), .B(new_n1121), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1116), .A2(KEYINPUT54), .A3(new_n1112), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT54), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT119), .B(G1996), .Z(new_n1132));
  OAI211_X1 g707(.A(new_n1014), .B(new_n1132), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n977), .A2(KEYINPUT118), .A3(new_n980), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT118), .B1(new_n977), .B2(new_n980), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT58), .B(G1341), .Z(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n631), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1142), .B(new_n631), .C1(new_n1133), .C2(new_n1137), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n577), .C2(new_n580), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT76), .B(G65), .Z(new_n1146));
  AOI22_X1  g721(.A1(new_n1146), .A2(new_n517), .B1(G78), .B2(G543), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n510), .B1(new_n1147), .B2(KEYINPUT77), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(new_n573), .B1(new_n603), .B2(G91), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n578), .B(KEYINPUT9), .ZN(new_n1150));
  OR2_X1    g725(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g726(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1956), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1088), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT56), .B(G2072), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1014), .B(new_n1157), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1154), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(KEYINPUT61), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1156), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n1159), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1138), .A2(KEYINPUT121), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1140), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1144), .A2(new_n1162), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT122), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1164), .A2(new_n1159), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1170), .A2(KEYINPUT61), .B1(new_n1140), .B2(new_n1166), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n1144), .A4(new_n1165), .ZN(new_n1173));
  AOI21_X1  g748(.A(G2067), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n758), .B2(new_n1031), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1175), .A2(KEYINPUT60), .A3(new_n622), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n622), .B1(new_n1175), .B2(KEYINPUT60), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1176), .A2(new_n1177), .B1(KEYINPUT60), .B2(new_n1175), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1169), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1175), .A2(new_n622), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1161), .B1(new_n1180), .B2(new_n1159), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1119), .A2(new_n1131), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1077), .A2(G286), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1124), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1120), .A2(G8), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1095), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1045), .A2(new_n1184), .A3(new_n1057), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1121), .A4(new_n1185), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1056), .A2(new_n1035), .A3(new_n591), .A4(new_n594), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1037), .B1(new_n1193), .B2(new_n1051), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1045), .A2(new_n1057), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1033), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1124), .A2(new_n1116), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1081), .A2(KEYINPUT62), .A3(new_n1083), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT62), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1192), .B(new_n1196), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1002), .B1(new_n1183), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n990), .B1(new_n987), .B2(new_n848), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n982), .B(KEYINPUT46), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT47), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n997), .B(KEYINPUT48), .Z(new_n1207));
  OAI21_X1  g782(.A(new_n1206), .B1(new_n995), .B2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n991), .A2(new_n811), .A3(new_n815), .A4(new_n818), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n986), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1208), .B1(new_n990), .B2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT127), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1202), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g788(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n1215), .B1(new_n896), .B2(new_n898), .ZN(new_n1216));
  NOR2_X1   g790(.A1(new_n962), .A2(new_n967), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1216), .A2(new_n1217), .ZN(G308));
  OR2_X1    g792(.A1(new_n1216), .A2(new_n1217), .ZN(G225));
endmodule


