//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT28), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT27), .B1(new_n206), .B2(KEYINPUT67), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G183gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n207), .B(new_n203), .C1(KEYINPUT67), .C2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n202), .A2(new_n213), .A3(KEYINPUT28), .A4(new_n203), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n218), .A2(KEYINPUT26), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(new_n206), .B2(new_n203), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n218), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G190gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n203), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n218), .B1(KEYINPUT23), .B2(new_n219), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n237), .B(new_n238), .C1(new_n229), .C2(new_n228), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n231), .A2(new_n236), .B1(new_n239), .B2(KEYINPUT25), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(G190gat), .A3(new_n232), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G190gat), .B2(new_n232), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  NOR4_X1   g042(.A1(new_n230), .A2(new_n242), .A3(new_n238), .A4(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n225), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G113gat), .A2(G120gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n246), .A2(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G127gat), .B(G134gat), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n252), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT25), .B1(new_n230), .B2(KEYINPUT66), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n236), .B(new_n237), .C1(new_n229), .C2(new_n228), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n231), .A2(KEYINPUT66), .A3(KEYINPUT25), .A4(new_n236), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n259), .A2(new_n260), .B1(new_n215), .B2(new_n224), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n252), .B(new_n254), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G227gat), .A2(G233gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT64), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT34), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT34), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n263), .A3(new_n266), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT33), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G15gat), .B(G43gat), .Z(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n274), .B(KEYINPUT32), .C1(new_n276), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT71), .A3(new_n272), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT36), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n269), .A3(new_n271), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT36), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n281), .A3(new_n283), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT37), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT22), .ZN(new_n296));
  INV_X1    g095(.A(G211gat), .ZN(new_n297));
  INV_X1    g096(.A(G218gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n295), .A3(new_n299), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT72), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(KEYINPUT72), .A3(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT74), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n245), .A2(new_n315), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT75), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n245), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n313), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n318), .A3(new_n308), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n294), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  OAI21_X1  g128(.A(KEYINPUT82), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT82), .ZN(new_n331));
  INV_X1    g130(.A(new_n329), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n261), .A2(new_n316), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n322), .B1(new_n321), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n333), .B1(new_n337), .B2(new_n313), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n331), .B(new_n332), .C1(new_n338), .C2(new_n294), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n294), .A3(new_n325), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT38), .ZN(new_n342));
  XOR2_X1   g141(.A(G1gat), .B(G29gat), .Z(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G141gat), .B(G148gat), .Z(new_n349));
  INV_X1    g148(.A(G155gat), .ZN(new_n350));
  INV_X1    g149(.A(G162gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT2), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G155gat), .B(G162gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n349), .A2(new_n354), .A3(new_n352), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT4), .B1(new_n255), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n357), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT3), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n262), .B(new_n365), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n255), .A2(new_n358), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n252), .A2(new_n254), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n252), .A2(new_n254), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n363), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n362), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n255), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n367), .A2(new_n378), .A3(new_n363), .A4(new_n379), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n368), .A2(new_n369), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n376), .A3(new_n369), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n348), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n369), .B1(new_n380), .B2(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n376), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n347), .A3(new_n382), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT6), .B(new_n348), .C1(new_n381), .C2(new_n383), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n335), .A2(new_n336), .A3(new_n312), .ZN(new_n394));
  INV_X1    g193(.A(new_n307), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(new_n305), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n321), .B2(new_n334), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT37), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n329), .A2(KEYINPUT38), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n399), .A2(new_n340), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n342), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT31), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G50gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n320), .B1(new_n364), .B2(new_n366), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n310), .A2(new_n311), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n303), .B2(new_n304), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n410), .A2(KEYINPUT3), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n411), .B2(new_n364), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n364), .B1(new_n410), .B2(new_n366), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n396), .A2(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n416), .A2(new_n417), .B1(G228gat), .B2(G233gat), .ZN(new_n418));
  OAI21_X1  g217(.A(G22gat), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n417), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n409), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n408), .A2(new_n412), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n406), .B1(new_n425), .B2(KEYINPUT80), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n406), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n427), .B(new_n430), .C1(new_n419), .C2(new_n424), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n312), .B1(new_n335), .B2(new_n336), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n332), .B1(new_n434), .B2(new_n333), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n392), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n338), .A2(new_n437), .A3(new_n329), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n361), .A2(new_n367), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n375), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(KEYINPUT39), .C1(new_n374), .C2(new_n375), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT39), .B1(new_n374), .B2(new_n375), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT81), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(new_n449), .A3(new_n375), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n347), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n441), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT40), .A3(new_n347), .A4(new_n450), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n452), .A2(new_n384), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n433), .B1(new_n440), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n293), .B1(new_n403), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n390), .A2(new_n391), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n433), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n431), .B1(new_n426), .B2(new_n428), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n284), .A3(new_n286), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT35), .B1(new_n462), .B2(new_n459), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n436), .A2(new_n438), .B1(new_n390), .B2(new_n391), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n288), .A2(new_n290), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n461), .A4(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n457), .A2(new_n460), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G29gat), .ZN(new_n469));
  INV_X1    g268(.A(G36gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT14), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(G29gat), .B2(G36gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G43gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G43gat), .ZN(new_n479));
  INV_X1    g278(.A(G50gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(KEYINPUT83), .A2(KEYINPUT15), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n483), .A2(new_n484), .B1(G43gat), .B2(G50gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G43gat), .A2(G50gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(G43gat), .A2(G50gat), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT15), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n475), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495));
  INV_X1    g294(.A(new_n489), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n484), .B1(new_n496), .B2(new_n487), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n483), .A2(new_n484), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n498), .A2(new_n487), .A3(new_n482), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n497), .B1(new_n499), .B2(new_n481), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n495), .B(new_n492), .C1(new_n500), .C2(new_n475), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n422), .A2(G15gat), .ZN(new_n504));
  INV_X1    g303(.A(G15gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G22gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(KEYINPUT16), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n510), .B2(G1gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(G8gat), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n509), .B(new_n512), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT17), .B1(new_n491), .B2(new_n493), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n519), .A3(new_n501), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n522), .A2(KEYINPUT18), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n485), .A2(new_n482), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n490), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n495), .B1(new_n531), .B2(new_n492), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n491), .A2(KEYINPUT85), .A3(new_n493), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n520), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n523), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n524), .B(KEYINPUT13), .Z(new_n536));
  AOI21_X1  g335(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  AOI211_X1 g337(.A(KEYINPUT90), .B(new_n538), .C1(new_n534), .C2(new_n523), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n525), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n503), .A2(new_n520), .A3(new_n521), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n524), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G197gat), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT11), .B(G169gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT91), .B1(new_n540), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n494), .A2(new_n519), .A3(new_n501), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n519), .B1(new_n494), .B2(new_n501), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n536), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n526), .A3(new_n536), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n550), .B1(new_n560), .B2(new_n541), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n559), .A2(new_n561), .A3(new_n562), .A4(new_n525), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(KEYINPUT89), .A3(new_n541), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n566), .A2(new_n559), .A3(new_n525), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n550), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT95), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G92gat), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G99gat), .ZN(new_n587));
  INV_X1    g386(.A(G106gat), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT8), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n581), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n581), .A2(new_n586), .A3(new_n591), .A4(new_n589), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n593), .A2(KEYINPUT96), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT96), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT97), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT8), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(G99gat), .B2(G106gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT95), .B(G92gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(new_n580), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n591), .B1(new_n603), .B2(new_n586), .ZN(new_n604));
  INV_X1    g403(.A(new_n594), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n593), .A2(KEYINPUT96), .A3(new_n594), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n598), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n597), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n503), .A2(new_n521), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT98), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(new_n598), .A3(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n503), .A2(new_n521), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n612), .A2(new_n533), .A3(new_n532), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n619), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n575), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n620), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n574), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(G71gat), .A2(G78gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G57gat), .B(G64gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G57gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G64gat), .ZN(new_n639));
  INV_X1    g438(.A(G64gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G57gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G71gat), .B(G78gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n636), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n519), .B1(KEYINPUT21), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n637), .A2(new_n645), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT21), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT20), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n649), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n659));
  XNOR2_X1  g458(.A(G183gat), .B(G211gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n631), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n646), .A2(KEYINPUT10), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n595), .A2(new_n596), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n646), .B1(new_n604), .B2(new_n605), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n593), .A2(new_n650), .A3(new_n594), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT10), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n666), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(new_n670), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n672), .B(new_n675), .C1(new_n676), .C2(new_n666), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  INV_X1    g477(.A(new_n666), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT10), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n593), .A2(new_n650), .A3(new_n594), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n650), .B1(new_n593), .B2(new_n594), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n646), .A4(new_n607), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n676), .A2(new_n666), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n678), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n677), .A2(new_n687), .ZN(new_n688));
  OR4_X1    g487(.A1(new_n468), .A2(new_n570), .A3(new_n665), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n458), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n508), .ZN(G1324gat));
  OAI21_X1  g490(.A(G8gat), .B1(new_n689), .B2(new_n439), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n689), .A2(new_n439), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT16), .B(G8gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT99), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n698));
  MUX2_X1   g497(.A(KEYINPUT100), .B(new_n698), .S(new_n696), .Z(new_n699));
  AOI22_X1  g498(.A1(new_n693), .A2(new_n697), .B1(new_n694), .B2(new_n699), .ZN(G1325gat));
  XOR2_X1   g499(.A(new_n292), .B(KEYINPUT101), .Z(new_n701));
  OAI21_X1  g500(.A(G15gat), .B1(new_n689), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n466), .A2(new_n505), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n689), .B2(new_n703), .ZN(G1326gat));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n461), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n570), .A2(new_n664), .A3(new_n688), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n468), .A2(new_n631), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n458), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n469), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT45), .Z(new_n714));
  NAND2_X1  g513(.A1(new_n463), .A2(new_n467), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n399), .A2(new_n340), .A3(new_n400), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(new_n391), .A3(new_n390), .A4(new_n392), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(KEYINPUT38), .B2(new_n341), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n455), .A2(new_n438), .A3(new_n436), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n461), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n292), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n459), .A2(KEYINPUT102), .A3(new_n433), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n464), .B2(new_n461), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n715), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT103), .B(new_n715), .C1(new_n721), .C2(new_n725), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n631), .A2(KEYINPUT44), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n468), .B2(new_n631), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n710), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n469), .B1(new_n733), .B2(new_n712), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n708), .B1(new_n714), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n734), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n713), .B(KEYINPUT45), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n711), .A2(new_n470), .A3(new_n440), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n731), .A2(new_n732), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n709), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT105), .B1(new_n744), .B2(new_n439), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G36gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n744), .A2(KEYINPUT105), .A3(new_n439), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n741), .B(new_n742), .C1(new_n746), .C2(new_n747), .ZN(G1329gat));
  NAND2_X1  g547(.A1(new_n477), .A2(new_n479), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n744), .B2(new_n292), .ZN(new_n750));
  INV_X1    g549(.A(new_n466), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n749), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n711), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n701), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n733), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n756), .A2(new_n749), .B1(new_n711), .B2(new_n752), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g557(.A1(new_n433), .A2(G50gat), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n711), .A2(new_n433), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n744), .A2(new_n759), .B1(G50gat), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g561(.A1(new_n728), .A2(new_n729), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n542), .A2(new_n543), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n557), .A2(new_n558), .B1(new_n764), .B2(KEYINPUT18), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n562), .B1(new_n765), .B2(new_n561), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n562), .A2(new_n559), .A3(new_n561), .A4(new_n525), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n569), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n688), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n665), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n458), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT106), .B(G57gat), .Z(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1332gat));
  INV_X1    g573(.A(new_n771), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n640), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n439), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n779), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT107), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n640), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n780), .A2(new_n777), .A3(new_n782), .A4(new_n640), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1333gat));
  INV_X1    g586(.A(G71gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n775), .A2(new_n788), .A3(new_n466), .ZN(new_n789));
  OAI21_X1  g588(.A(G71gat), .B1(new_n771), .B2(new_n701), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(KEYINPUT50), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n433), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n722), .A2(new_n724), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n457), .A2(new_n799), .B1(new_n463), .B2(new_n467), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(new_n631), .ZN(new_n801));
  INV_X1    g600(.A(new_n631), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n726), .A2(KEYINPUT109), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n664), .A2(new_n768), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n801), .A2(new_n803), .A3(new_n808), .A4(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n580), .A3(new_n712), .A4(new_n688), .ZN(new_n811));
  INV_X1    g610(.A(new_n664), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n570), .A3(new_n688), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT108), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n731), .B2(new_n732), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G85gat), .B1(new_n817), .B2(new_n458), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n818), .ZN(G1336gat));
  NOR2_X1   g618(.A1(new_n439), .A2(new_n769), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n576), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n807), .B2(new_n809), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n602), .B1(new_n816), .B2(new_n440), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n822), .B2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1337gat));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n587), .A3(new_n466), .A4(new_n688), .ZN(new_n829));
  OAI21_X1  g628(.A(G99gat), .B1(new_n817), .B2(new_n701), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1338gat));
  NOR3_X1   g630(.A1(new_n461), .A2(G106gat), .A3(new_n769), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n810), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT111), .B(G106gat), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n461), .B(new_n815), .C1(new_n731), .C2(new_n732), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(KEYINPUT112), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n433), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n836), .A2(new_n834), .ZN(new_n840));
  INV_X1    g639(.A(new_n832), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n807), .B2(new_n809), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(G1339gat));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n554), .A2(new_n555), .A3(new_n536), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n548), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n688), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n845), .B1(new_n564), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT114), .B(new_n849), .C1(new_n553), .C2(new_n563), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n675), .B1(new_n685), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n683), .A2(new_n684), .A3(new_n679), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n672), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT55), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT113), .A3(new_n677), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n857), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT113), .B1(new_n858), .B2(new_n677), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n768), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n802), .B1(new_n853), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n848), .B1(new_n766), .B2(new_n767), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n858), .A2(new_n677), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n859), .A3(new_n862), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n631), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n812), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  AND4_X1   g673(.A1(new_n570), .A2(new_n664), .A3(new_n631), .A4(new_n769), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n433), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n877), .A2(new_n712), .A3(new_n439), .A4(new_n466), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n570), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT115), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n458), .B1(new_n874), .B2(new_n876), .ZN(new_n881));
  INV_X1    g680(.A(new_n462), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n439), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n768), .A2(new_n248), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(G1340gat));
  OAI21_X1  g685(.A(G120gat), .B1(new_n878), .B2(new_n769), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n688), .A2(new_n249), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT116), .ZN(G1341gat));
  OAI21_X1  g689(.A(G127gat), .B1(new_n878), .B2(new_n812), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n812), .A2(G127gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n884), .B2(new_n892), .ZN(G1342gat));
  INV_X1    g692(.A(G134gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n802), .A2(new_n439), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT117), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n883), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT118), .ZN(new_n900));
  OAI21_X1  g699(.A(G134gat), .B1(new_n878), .B2(new_n631), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n900), .B(new_n901), .C1(KEYINPUT56), .C2(new_n898), .ZN(G1343gat));
  INV_X1    g701(.A(G141gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n292), .A2(new_n712), .A3(new_n439), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n862), .A2(new_n677), .A3(new_n858), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n564), .B2(new_n569), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n849), .B1(new_n553), .B2(new_n563), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n631), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n848), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n553), .B2(new_n563), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n865), .A2(new_n630), .A3(new_n910), .A4(new_n626), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n664), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT57), .B(new_n433), .C1(new_n912), .C2(new_n875), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n850), .B1(new_n766), .B2(new_n767), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT114), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n907), .A2(new_n845), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n866), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n873), .B1(new_n918), .B2(new_n631), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n876), .B1(new_n919), .B2(new_n664), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT57), .B1(new_n920), .B2(new_n433), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n914), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n461), .B1(new_n874), .B2(new_n876), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT119), .B1(new_n924), .B2(KEYINPUT57), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n904), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n903), .B1(new_n926), .B2(new_n768), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n755), .A2(new_n461), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(new_n439), .A3(new_n881), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(new_n903), .A3(new_n768), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n927), .A2(KEYINPUT58), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT58), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1344gat));
  INV_X1    g732(.A(G148gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n934), .A3(new_n688), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G148gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n926), .B2(new_n688), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n904), .A2(new_n769), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT57), .ZN(new_n940));
  INV_X1    g739(.A(new_n905), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n907), .B1(new_n768), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n911), .B1(new_n942), .B2(new_n802), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n875), .B1(new_n943), .B2(new_n812), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n944), .B2(new_n461), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n924), .A2(KEYINPUT57), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND4_X1   g746(.A1(new_n946), .A2(new_n920), .A3(KEYINPUT57), .A4(new_n433), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n939), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n936), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n935), .B1(new_n938), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT121), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(new_n935), .C1(new_n938), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1345gat));
  NAND3_X1  g754(.A1(new_n929), .A2(new_n350), .A3(new_n664), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n926), .A2(new_n664), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n350), .ZN(G1346gat));
  NAND4_X1  g757(.A1(new_n928), .A2(new_n351), .A3(new_n881), .A4(new_n897), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n926), .A2(new_n802), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n351), .ZN(G1347gat));
  NAND2_X1  g760(.A1(new_n440), .A2(new_n458), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(new_n751), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT124), .Z(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n877), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(new_n216), .A3(new_n570), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n712), .B1(new_n874), .B2(new_n876), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n882), .A2(new_n440), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT122), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n967), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n768), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n966), .B1(new_n976), .B2(new_n216), .ZN(G1348gat));
  OAI21_X1  g776(.A(G176gat), .B1(new_n965), .B2(new_n769), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n688), .A2(new_n217), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n974), .B2(new_n979), .ZN(G1349gat));
  OAI21_X1  g779(.A(G183gat), .B1(new_n965), .B2(new_n812), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n664), .A2(new_n202), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n970), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g783(.A1(new_n975), .A2(new_n203), .A3(new_n802), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n964), .A2(new_n877), .A3(new_n802), .ZN(new_n986));
  XNOR2_X1  g785(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n986), .A2(G190gat), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n986), .B2(G190gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n985), .B(new_n992), .C1(new_n989), .C2(new_n988), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1351gat));
  AND2_X1   g793(.A1(new_n928), .A2(new_n967), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n995), .A2(new_n440), .ZN(new_n996));
  AOI21_X1  g795(.A(G197gat), .B1(new_n996), .B2(new_n768), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n947), .A2(new_n948), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n755), .A2(new_n962), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n768), .A2(G197gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(G1352gat));
  INV_X1    g802(.A(G204gat), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n995), .A2(new_n1004), .A3(new_n820), .ZN(new_n1005));
  XOR2_X1   g804(.A(new_n1005), .B(KEYINPUT62), .Z(new_n1006));
  OAI21_X1  g805(.A(G204gat), .B1(new_n1000), .B2(new_n769), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1353gat));
  NAND3_X1  g807(.A1(new_n996), .A2(new_n297), .A3(new_n664), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n998), .A2(new_n664), .A3(new_n999), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1010), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT63), .B1(new_n1010), .B2(G211gat), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(G1354gat));
  OAI21_X1  g812(.A(G218gat), .B1(new_n1000), .B2(new_n631), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n298), .A3(new_n802), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(G1355gat));
endmodule


