

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X2 U553 ( .A1(n525), .A2(G2104), .ZN(n888) );
  NOR2_X1 U554 ( .A1(n529), .A2(n528), .ZN(G160) );
  XNOR2_X1 U555 ( .A(n531), .B(KEYINPUT0), .ZN(n663) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n647) );
  XNOR2_X1 U557 ( .A(KEYINPUT91), .B(n812), .ZN(n520) );
  OR2_X1 U558 ( .A1(n698), .A2(n699), .ZN(n701) );
  NOR2_X1 U559 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U560 ( .A1(n790), .A2(n693), .ZN(n699) );
  BUF_X1 U561 ( .A(n699), .Z(n739) );
  OR2_X1 U562 ( .A1(n663), .A2(n535), .ZN(n536) );
  NAND2_X1 U563 ( .A1(n520), .A2(n813), .ZN(n814) );
  INV_X1 U564 ( .A(G543), .ZN(n531) );
  INV_X1 U565 ( .A(n536), .ZN(n650) );
  NOR2_X1 U566 ( .A1(n541), .A2(n540), .ZN(G171) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n521), .Z(n887) );
  NAND2_X1 U569 ( .A1(n887), .A2(G137), .ZN(n524) );
  INV_X1 U570 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U571 ( .A1(G101), .A2(n888), .ZN(n522) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n529) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n525), .ZN(n893) );
  NAND2_X1 U575 ( .A1(G125), .A2(n893), .ZN(n527) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U577 ( .A1(G113), .A2(n891), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  INV_X1 U579 ( .A(G651), .ZN(n535) );
  NOR2_X1 U580 ( .A1(G543), .A2(n535), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n530), .Z(n662) );
  NAND2_X1 U582 ( .A1(G64), .A2(n662), .ZN(n534) );
  NOR2_X1 U583 ( .A1(G651), .A2(n663), .ZN(n532) );
  XNOR2_X1 U584 ( .A(KEYINPUT64), .B(n532), .ZN(n656) );
  NAND2_X1 U585 ( .A1(G52), .A2(n656), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U587 ( .A1(G90), .A2(n647), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G77), .A2(n650), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U590 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  XOR2_X1 U591 ( .A(G2443), .B(G2446), .Z(n543) );
  XNOR2_X1 U592 ( .A(G2427), .B(G2451), .ZN(n542) );
  XNOR2_X1 U593 ( .A(n543), .B(n542), .ZN(n549) );
  XOR2_X1 U594 ( .A(G2430), .B(G2454), .Z(n545) );
  XNOR2_X1 U595 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U596 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U597 ( .A(G2435), .B(G2438), .Z(n546) );
  XNOR2_X1 U598 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U599 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U600 ( .A1(G14), .A2(n550), .ZN(G401) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  NAND2_X1 U603 ( .A1(n887), .A2(G138), .ZN(n556) );
  NAND2_X1 U604 ( .A1(G114), .A2(n891), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G102), .A2(n888), .ZN(n551) );
  AND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G126), .A2(n893), .ZN(n553) );
  AND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U610 ( .A(n557), .B(KEYINPUT85), .ZN(G164) );
  NAND2_X1 U611 ( .A1(G65), .A2(n662), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G53), .A2(n656), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U614 ( .A(KEYINPUT65), .B(n560), .ZN(n564) );
  NAND2_X1 U615 ( .A1(G91), .A2(n647), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G78), .A2(n650), .ZN(n561) );
  AND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U620 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n832) );
  NAND2_X1 U622 ( .A1(n832), .A2(G567), .ZN(n566) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U624 ( .A1(n647), .A2(G81), .ZN(n567) );
  XNOR2_X1 U625 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G68), .A2(n650), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n571) );
  XOR2_X1 U628 ( .A(KEYINPUT66), .B(KEYINPUT13), .Z(n570) );
  XNOR2_X1 U629 ( .A(n571), .B(n570), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n662), .A2(G56), .ZN(n572) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G43), .A2(n656), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n920) );
  INV_X1 U635 ( .A(G860), .ZN(n605) );
  OR2_X1 U636 ( .A1(n920), .A2(n605), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G868), .A2(G171), .ZN(n587) );
  NAND2_X1 U638 ( .A1(n650), .A2(G79), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT67), .B(n577), .Z(n579) );
  NAND2_X1 U640 ( .A1(G54), .A2(n656), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT68), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G92), .A2(n647), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G66), .A2(n662), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X2 U647 ( .A(KEYINPUT15), .B(n585), .Z(n933) );
  INV_X1 U648 ( .A(G868), .ZN(n609) );
  NAND2_X1 U649 ( .A1(n933), .A2(n609), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U651 ( .A(n588), .B(KEYINPUT69), .ZN(G284) );
  NAND2_X1 U652 ( .A1(n662), .A2(G63), .ZN(n589) );
  XNOR2_X1 U653 ( .A(KEYINPUT71), .B(n589), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G51), .A2(n656), .ZN(n590) );
  XOR2_X1 U655 ( .A(n590), .B(KEYINPUT72), .Z(n591) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT6), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(KEYINPUT73), .ZN(n601) );
  NAND2_X1 U659 ( .A1(G89), .A2(n647), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n595), .B(KEYINPUT70), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n596), .B(KEYINPUT4), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G76), .A2(n650), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U664 ( .A(KEYINPUT5), .B(n599), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U666 ( .A(n602), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U667 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U668 ( .A1(G286), .A2(n609), .ZN(n604) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U670 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U671 ( .A1(G559), .A2(n605), .ZN(n606) );
  XNOR2_X1 U672 ( .A(KEYINPUT74), .B(n606), .ZN(n607) );
  NAND2_X1 U673 ( .A1(n607), .A2(n933), .ZN(n608) );
  XNOR2_X1 U674 ( .A(KEYINPUT16), .B(n608), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G559), .A2(n609), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n933), .A2(n610), .ZN(n611) );
  XNOR2_X1 U677 ( .A(n611), .B(KEYINPUT75), .ZN(n613) );
  NOR2_X1 U678 ( .A1(n920), .A2(G868), .ZN(n612) );
  NOR2_X1 U679 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U680 ( .A1(n893), .A2(G123), .ZN(n614) );
  XNOR2_X1 U681 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G111), .A2(n891), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U684 ( .A1(G135), .A2(n887), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G99), .A2(n888), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n996) );
  XNOR2_X1 U688 ( .A(n996), .B(G2096), .ZN(n622) );
  INV_X1 U689 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U691 ( .A1(n933), .A2(G559), .ZN(n672) );
  XNOR2_X1 U692 ( .A(n920), .B(n672), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n623), .A2(G860), .ZN(n630) );
  NAND2_X1 U694 ( .A1(G93), .A2(n647), .ZN(n625) );
  NAND2_X1 U695 ( .A1(G80), .A2(n650), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G67), .A2(n662), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G55), .A2(n656), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n674) );
  XNOR2_X1 U701 ( .A(n630), .B(n674), .ZN(G145) );
  AND2_X1 U702 ( .A1(n662), .A2(G60), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G85), .A2(n647), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G72), .A2(n650), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U707 ( .A1(G47), .A2(n656), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U709 ( .A1(G73), .A2(n650), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT2), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n638), .B(KEYINPUT78), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G86), .A2(n647), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U714 ( .A1(G61), .A2(n662), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G48), .A2(n656), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U718 ( .A(KEYINPUT79), .B(n645), .ZN(G305) );
  NAND2_X1 U719 ( .A1(n656), .A2(G50), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT80), .ZN(n655) );
  NAND2_X1 U721 ( .A1(G88), .A2(n647), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G62), .A2(n662), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U724 ( .A1(G75), .A2(n650), .ZN(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT81), .B(n651), .ZN(n652) );
  NOR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(G303) );
  INV_X1 U728 ( .A(G303), .ZN(G166) );
  NAND2_X1 U729 ( .A1(n656), .A2(G49), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(KEYINPUT76), .ZN(n660) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n658) );
  XOR2_X1 U732 ( .A(KEYINPUT77), .B(n658), .Z(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n663), .A2(G87), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(G288) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(G290), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(G305), .ZN(n669) );
  XNOR2_X1 U739 ( .A(G166), .B(G299), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n667), .B(G288), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n920), .B(n674), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n902) );
  XOR2_X1 U744 ( .A(n902), .B(n672), .Z(n673) );
  NAND2_X1 U745 ( .A1(G868), .A2(n673), .ZN(n676) );
  OR2_X1 U746 ( .A1(n674), .A2(G868), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n681) );
  NOR2_X1 U755 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U756 ( .A1(G108), .A2(n682), .ZN(n837) );
  NAND2_X1 U757 ( .A1(G567), .A2(n837), .ZN(n689) );
  NAND2_X1 U758 ( .A1(G132), .A2(G82), .ZN(n683) );
  XNOR2_X1 U759 ( .A(n683), .B(KEYINPUT82), .ZN(n684) );
  XNOR2_X1 U760 ( .A(n684), .B(KEYINPUT22), .ZN(n685) );
  NOR2_X1 U761 ( .A1(G218), .A2(n685), .ZN(n686) );
  XOR2_X1 U762 ( .A(KEYINPUT83), .B(n686), .Z(n687) );
  NAND2_X1 U763 ( .A1(G96), .A2(n687), .ZN(n838) );
  NAND2_X1 U764 ( .A1(G2106), .A2(n838), .ZN(n688) );
  NAND2_X1 U765 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U766 ( .A(KEYINPUT84), .B(n690), .Z(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n692) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U769 ( .A1(n692), .A2(n691), .ZN(n836) );
  NAND2_X1 U770 ( .A1(n836), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n790) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n791) );
  INV_X1 U773 ( .A(n791), .ZN(n693) );
  NAND2_X1 U774 ( .A1(G8), .A2(n739), .ZN(n775) );
  INV_X1 U775 ( .A(n699), .ZN(n703) );
  NAND2_X1 U776 ( .A1(n703), .A2(G2072), .ZN(n694) );
  XOR2_X1 U777 ( .A(KEYINPUT27), .B(n694), .Z(n716) );
  NAND2_X1 U778 ( .A1(G1956), .A2(n739), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n716), .A2(n714), .ZN(n695) );
  NAND2_X1 U780 ( .A1(n695), .A2(G299), .ZN(n696) );
  XNOR2_X1 U781 ( .A(n696), .B(KEYINPUT93), .ZN(n697) );
  XNOR2_X1 U782 ( .A(KEYINPUT28), .B(n697), .ZN(n723) );
  INV_X1 U783 ( .A(G2067), .ZN(n698) );
  NAND2_X1 U784 ( .A1(G1348), .A2(n699), .ZN(n700) );
  NAND2_X1 U785 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U786 ( .A(KEYINPUT94), .B(n702), .Z(n710) );
  OR2_X1 U787 ( .A1(n933), .A2(n710), .ZN(n709) );
  AND2_X1 U788 ( .A1(n703), .A2(G1996), .ZN(n704) );
  XOR2_X1 U789 ( .A(n704), .B(KEYINPUT26), .Z(n706) );
  NAND2_X1 U790 ( .A1(n739), .A2(G1341), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U792 ( .A1(n920), .A2(n707), .ZN(n708) );
  NAND2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n710), .A2(n933), .ZN(n711) );
  NAND2_X1 U795 ( .A1(n712), .A2(n711), .ZN(n720) );
  INV_X1 U796 ( .A(KEYINPUT95), .ZN(n718) );
  INV_X1 U797 ( .A(G299), .ZN(n713) );
  AND2_X1 U798 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U799 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U800 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U801 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U802 ( .A(KEYINPUT96), .B(n721), .ZN(n722) );
  XNOR2_X1 U803 ( .A(n724), .B(KEYINPUT29), .ZN(n729) );
  NOR2_X1 U804 ( .A1(n703), .A2(G1961), .ZN(n725) );
  XOR2_X1 U805 ( .A(KEYINPUT92), .B(n725), .Z(n727) );
  XNOR2_X1 U806 ( .A(KEYINPUT25), .B(G2078), .ZN(n979) );
  NAND2_X1 U807 ( .A1(n703), .A2(n979), .ZN(n726) );
  NAND2_X1 U808 ( .A1(n727), .A2(n726), .ZN(n733) );
  NAND2_X1 U809 ( .A1(G171), .A2(n733), .ZN(n728) );
  NAND2_X1 U810 ( .A1(n729), .A2(n728), .ZN(n738) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n775), .ZN(n750) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n739), .ZN(n747) );
  NOR2_X1 U813 ( .A1(n750), .A2(n747), .ZN(n730) );
  NAND2_X1 U814 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  NOR2_X1 U816 ( .A1(G168), .A2(n732), .ZN(n735) );
  NOR2_X1 U817 ( .A1(G171), .A2(n733), .ZN(n734) );
  NOR2_X1 U818 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(n736), .Z(n737) );
  NAND2_X1 U820 ( .A1(n738), .A2(n737), .ZN(n748) );
  NAND2_X1 U821 ( .A1(G286), .A2(n748), .ZN(n744) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n775), .ZN(n741) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U824 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U825 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U826 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U827 ( .A1(n745), .A2(G8), .ZN(n746) );
  XNOR2_X1 U828 ( .A(n746), .B(KEYINPUT32), .ZN(n767) );
  NAND2_X1 U829 ( .A1(G8), .A2(n747), .ZN(n752) );
  INV_X1 U830 ( .A(n748), .ZN(n749) );
  NAND2_X1 U831 ( .A1(n752), .A2(n751), .ZN(n768) );
  NAND2_X1 U832 ( .A1(G288), .A2(G1976), .ZN(n753) );
  XOR2_X1 U833 ( .A(KEYINPUT98), .B(n753), .Z(n928) );
  INV_X1 U834 ( .A(n928), .ZN(n754) );
  AND2_X1 U835 ( .A1(n768), .A2(n754), .ZN(n755) );
  NAND2_X1 U836 ( .A1(n767), .A2(n755), .ZN(n759) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n917) );
  XOR2_X1 U838 ( .A(KEYINPUT97), .B(n917), .Z(n756) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n929) );
  NOR2_X1 U840 ( .A1(n756), .A2(n929), .ZN(n757) );
  OR2_X1 U841 ( .A1(n928), .A2(n757), .ZN(n758) );
  NAND2_X1 U842 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U843 ( .A(n760), .B(KEYINPUT99), .ZN(n761) );
  NOR2_X1 U844 ( .A1(n775), .A2(n761), .ZN(n762) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n762), .ZN(n765) );
  NAND2_X1 U846 ( .A1(n929), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U847 ( .A1(n763), .A2(n775), .ZN(n764) );
  NOR2_X1 U848 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n912) );
  AND2_X1 U850 ( .A1(n766), .A2(n912), .ZN(n779) );
  NAND2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n771) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U853 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n772), .A2(n775), .ZN(n777) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XOR2_X1 U857 ( .A(n773), .B(KEYINPUT24), .Z(n774) );
  OR2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U859 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U860 ( .A1(n779), .A2(n778), .ZN(n815) );
  XNOR2_X1 U861 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NAND2_X1 U862 ( .A1(G140), .A2(n887), .ZN(n781) );
  NAND2_X1 U863 ( .A1(G104), .A2(n888), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U866 ( .A1(G128), .A2(n893), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G116), .A2(n891), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U869 ( .A(n785), .B(KEYINPUT35), .Z(n786) );
  NOR2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U871 ( .A(KEYINPUT36), .B(n788), .Z(n789) );
  XNOR2_X1 U872 ( .A(KEYINPUT87), .B(n789), .ZN(n883) );
  NOR2_X1 U873 ( .A1(n825), .A2(n883), .ZN(n1002) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U875 ( .A(n792), .B(KEYINPUT86), .Z(n810) );
  INV_X1 U876 ( .A(n810), .ZN(n827) );
  NAND2_X1 U877 ( .A1(n1002), .A2(n827), .ZN(n823) );
  XNOR2_X1 U878 ( .A(KEYINPUT88), .B(G1991), .ZN(n970) );
  NAND2_X1 U879 ( .A1(G119), .A2(n893), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G131), .A2(n887), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G107), .A2(n891), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G95), .A2(n888), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n866) );
  AND2_X1 U886 ( .A1(n970), .A2(n866), .ZN(n809) );
  NAND2_X1 U887 ( .A1(G105), .A2(n888), .ZN(n799) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  XNOR2_X1 U889 ( .A(n800), .B(KEYINPUT89), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G129), .A2(n893), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U892 ( .A1(G141), .A2(n887), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G117), .A2(n891), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U896 ( .A(KEYINPUT90), .B(n807), .Z(n867) );
  AND2_X1 U897 ( .A1(n867), .A2(G1996), .ZN(n808) );
  NOR2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n994) );
  NOR2_X1 U899 ( .A1(n810), .A2(n994), .ZN(n819) );
  INV_X1 U900 ( .A(n819), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n823), .A2(n811), .ZN(n812) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n916) );
  NAND2_X1 U903 ( .A1(n916), .A2(n827), .ZN(n813) );
  OR2_X2 U904 ( .A1(n815), .A2(n814), .ZN(n830) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U906 ( .A1(n970), .A2(n866), .ZN(n997) );
  NOR2_X1 U907 ( .A1(n816), .A2(n997), .ZN(n817) );
  XOR2_X1 U908 ( .A(KEYINPUT101), .B(n817), .Z(n818) );
  NOR2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n821) );
  NOR2_X1 U910 ( .A1(n867), .A2(G1996), .ZN(n820) );
  XNOR2_X1 U911 ( .A(n820), .B(KEYINPUT100), .ZN(n991) );
  NOR2_X1 U912 ( .A1(n821), .A2(n991), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U915 ( .A1(n825), .A2(n883), .ZN(n1005) );
  NAND2_X1 U916 ( .A1(n826), .A2(n1005), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U919 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(n832), .A2(G2106), .ZN(n833) );
  XNOR2_X1 U921 ( .A(n833), .B(KEYINPUT102), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U923 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U927 ( .A(G132), .ZN(G219) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n839), .B(KEYINPUT103), .ZN(G261) );
  INV_X1 U934 ( .A(G261), .ZN(G325) );
  XOR2_X1 U935 ( .A(KEYINPUT41), .B(G1956), .Z(n841) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U938 ( .A(n842), .B(KEYINPUT105), .Z(n844) );
  XNOR2_X1 U939 ( .A(G1961), .B(G1971), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U941 ( .A(G1976), .B(G1981), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1966), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U945 ( .A(KEYINPUT104), .B(G2474), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n852) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(G227) );
  NAND2_X1 U956 ( .A1(n893), .A2(G124), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G112), .A2(n891), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U960 ( .A1(G136), .A2(n887), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G100), .A2(n888), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U963 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n869) );
  XOR2_X1 U965 ( .A(n867), .B(n866), .Z(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n882) );
  XNOR2_X1 U967 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G142), .A2(n887), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G106), .A2(n888), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT45), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G130), .A2(n893), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G118), .A2(n891), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U976 ( .A(KEYINPUT106), .B(n877), .ZN(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U978 ( .A(G160), .B(n880), .Z(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n883), .B(n996), .ZN(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U982 ( .A(n886), .B(G162), .Z(n900) );
  NAND2_X1 U983 ( .A1(G139), .A2(n887), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U986 ( .A1(n891), .A2(G115), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT109), .B(n892), .Z(n895) );
  NAND2_X1 U988 ( .A1(n893), .A2(G127), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n1009) );
  XNOR2_X1 U992 ( .A(G164), .B(n1009), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U994 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n933), .B(G286), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U997 ( .A(n904), .B(G171), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n906) );
  XOR2_X1 U1000 ( .A(KEYINPUT49), .B(n906), .Z(n907) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n907), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n908), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n909), .B(KEYINPUT110), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G171), .ZN(G301) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1009 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1027) );
  XNOR2_X1 U1010 ( .A(KEYINPUT56), .B(G16), .ZN(n941) );
  XNOR2_X1 U1011 ( .A(G1966), .B(G168), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(KEYINPUT120), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(KEYINPUT57), .B(n915), .ZN(n938) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(G171), .B(G1961), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(G1971), .A2(G303), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(G1341), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G1956), .B(G299), .Z(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT121), .B(n925), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n930), .B(KEYINPUT122), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n936) );
  INV_X1 U1028 ( .A(n933), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G1348), .B(n934), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1032 ( .A(KEYINPUT123), .B(n939), .Z(n940) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n1025) );
  XOR2_X1 U1034 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n964) );
  XNOR2_X1 U1035 ( .A(G1341), .B(G19), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(G1981), .B(G6), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT124), .B(n944), .Z(n946) );
  XNOR2_X1 U1039 ( .A(G1956), .B(G20), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n950) );
  XOR2_X1 U1041 ( .A(KEYINPUT125), .B(G4), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(n951), .B(KEYINPUT60), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G22), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G23), .B(G1976), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1049 ( .A(G1986), .B(G24), .Z(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT58), .B(n956), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G21), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G5), .B(G1961), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n964), .B(n963), .ZN(n966) );
  INV_X1 U1058 ( .A(G16), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n967), .ZN(n1023) );
  XOR2_X1 U1061 ( .A(G34), .B(KEYINPUT118), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G2084), .B(KEYINPUT54), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n986) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n984) );
  XOR2_X1 U1065 ( .A(n970), .B(G25), .Z(n978) );
  XNOR2_X1 U1066 ( .A(G2067), .B(G26), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G33), .B(G2072), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(G28), .A2(n973), .ZN(n976) );
  XOR2_X1 U1070 ( .A(KEYINPUT117), .B(G1996), .Z(n974) );
  XNOR2_X1 U1071 ( .A(G32), .B(n974), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1074 ( .A(G27), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT55), .B(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n988), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n989), .B(KEYINPUT119), .ZN(n1021) );
  XOR2_X1 U1082 ( .A(G2090), .B(G162), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(KEYINPUT113), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT51), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1007) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT111), .B(n998), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(G160), .B(G2084), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT112), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(KEYINPUT114), .B(n1008), .ZN(n1014) );
  XOR2_X1 U1096 ( .A(G2072), .B(n1009), .Z(n1011) );
  XOR2_X1 U1097 ( .A(G164), .B(G2078), .Z(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(n1015), .B(KEYINPUT115), .Z(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1017), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT116), .B(n1018), .Z(n1019) );
  NAND2_X1 U1105 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(n1027), .B(n1026), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

