

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770;

  NAND2_X1 U369 ( .A1(n416), .A2(n415), .ZN(n553) );
  NOR2_X2 U370 ( .A1(n694), .A2(n587), .ZN(n588) );
  NOR2_X1 U371 ( .A1(n539), .A2(n379), .ZN(n405) );
  XNOR2_X1 U372 ( .A(n594), .B(n434), .ZN(n701) );
  BUF_X1 U373 ( .A(G104), .Z(n347) );
  XNOR2_X1 U374 ( .A(n752), .B(n428), .ZN(n483) );
  XNOR2_X1 U375 ( .A(n472), .B(n471), .ZN(n751) );
  NAND2_X1 U376 ( .A1(n729), .A2(G472), .ZN(n664) );
  AND2_X2 U377 ( .A1(n638), .A2(n639), .ZN(n729) );
  XNOR2_X1 U378 ( .A(G140), .B(n347), .ZN(n514) );
  AND2_X2 U379 ( .A1(n655), .A2(n652), .ZN(n561) );
  NOR2_X2 U380 ( .A1(n647), .A2(n742), .ZN(n648) );
  NOR2_X2 U381 ( .A1(n665), .A2(n742), .ZN(n667) );
  NOR2_X2 U382 ( .A1(n659), .A2(n742), .ZN(n661) );
  XNOR2_X2 U383 ( .A(G113), .B(G119), .ZN(n418) );
  OR2_X2 U384 ( .A1(n701), .A2(n700), .ZN(n539) );
  XNOR2_X1 U385 ( .A(G953), .B(KEYINPUT64), .ZN(n349) );
  XNOR2_X1 U386 ( .A(n412), .B(n411), .ZN(n373) );
  XNOR2_X1 U387 ( .A(n543), .B(KEYINPUT31), .ZN(n681) );
  NOR2_X1 U388 ( .A1(n626), .A2(n675), .ZN(n586) );
  AND2_X1 U389 ( .A1(n388), .A2(n386), .ZN(n385) );
  XNOR2_X1 U390 ( .A(n420), .B(n419), .ZN(n472) );
  INV_X2 U391 ( .A(n349), .ZN(n440) );
  INV_X2 U392 ( .A(G128), .ZN(n406) );
  BUF_X1 U393 ( .A(n533), .Z(n348) );
  XNOR2_X1 U394 ( .A(n553), .B(KEYINPUT105), .ZN(n533) );
  INV_X2 U395 ( .A(G125), .ZN(n380) );
  NAND2_X1 U396 ( .A1(n348), .A2(n532), .ZN(n350) );
  NAND2_X1 U397 ( .A1(n533), .A2(n532), .ZN(n655) );
  BUF_X1 U398 ( .A(n729), .Z(n738) );
  INV_X1 U399 ( .A(KEYINPUT83), .ZN(n369) );
  INV_X1 U400 ( .A(KEYINPUT22), .ZN(n417) );
  NAND2_X1 U401 ( .A1(n695), .A2(KEYINPUT103), .ZN(n391) );
  AND2_X1 U402 ( .A1(n552), .A2(n399), .ZN(n396) );
  XNOR2_X1 U403 ( .A(KEYINPUT74), .B(KEYINPUT100), .ZN(n458) );
  XNOR2_X1 U404 ( .A(n374), .B(n376), .ZN(n464) );
  XNOR2_X1 U405 ( .A(n423), .B(G146), .ZN(n376) );
  XNOR2_X1 U406 ( .A(n375), .B(n457), .ZN(n374) );
  XNOR2_X1 U407 ( .A(n503), .B(n351), .ZN(n467) );
  AND2_X1 U408 ( .A1(n685), .A2(n359), .ZN(n413) );
  AND2_X1 U409 ( .A1(n368), .A2(n686), .ZN(n367) );
  XNOR2_X1 U410 ( .A(n467), .B(n442), .ZN(n759) );
  XNOR2_X1 U411 ( .A(n421), .B(G116), .ZN(n419) );
  INV_X1 U412 ( .A(KEYINPUT69), .ZN(n421) );
  AND2_X1 U413 ( .A1(n691), .A2(n410), .ZN(n409) );
  XNOR2_X1 U414 ( .A(n407), .B(n576), .ZN(n609) );
  NAND2_X1 U415 ( .A1(n575), .A2(n692), .ZN(n407) );
  XNOR2_X1 U416 ( .A(n426), .B(n425), .ZN(n752) );
  XNOR2_X1 U417 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U418 ( .A(G119), .B(G128), .ZN(n443) );
  XNOR2_X1 U419 ( .A(n588), .B(KEYINPUT41), .ZN(n721) );
  NAND2_X2 U420 ( .A1(n385), .A2(n381), .ZN(n604) );
  NAND2_X1 U421 ( .A1(n384), .A2(n382), .ZN(n381) );
  NOR2_X1 U422 ( .A1(n596), .A2(n595), .ZN(n619) );
  NAND2_X1 U423 ( .A1(n662), .A2(n486), .ZN(n469) );
  INV_X1 U424 ( .A(n623), .ZN(n415) );
  AND2_X1 U425 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U426 ( .A1(n392), .A2(n390), .ZN(n389) );
  NOR2_X1 U427 ( .A1(G953), .A2(G237), .ZN(n518) );
  INV_X1 U428 ( .A(G237), .ZN(n485) );
  XOR2_X1 U429 ( .A(G122), .B(G143), .Z(n513) );
  NAND2_X1 U430 ( .A1(G234), .A2(G237), .ZN(n492) );
  INV_X1 U431 ( .A(KEYINPUT85), .ZN(n383) );
  NAND2_X1 U432 ( .A1(n387), .A2(KEYINPUT85), .ZN(n386) );
  INV_X1 U433 ( .A(n692), .ZN(n387) );
  NOR2_X1 U434 ( .A1(G902), .A2(n735), .ZN(n529) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n662) );
  NAND2_X1 U436 ( .A1(n466), .A2(n465), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n467), .B(n472), .ZN(n377) );
  NAND2_X2 U438 ( .A1(n366), .A2(n364), .ZN(n765) );
  NAND2_X1 U439 ( .A1(n365), .A2(n369), .ZN(n364) );
  AND2_X1 U440 ( .A1(n370), .A2(n367), .ZN(n366) );
  XNOR2_X1 U441 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U442 ( .A(n474), .B(G134), .ZN(n503) );
  XNOR2_X1 U443 ( .A(n431), .B(n759), .ZN(n730) );
  XOR2_X1 U444 ( .A(KEYINPUT77), .B(KEYINPUT18), .Z(n475) );
  XNOR2_X1 U445 ( .A(n405), .B(KEYINPUT33), .ZN(n720) );
  XNOR2_X1 U446 ( .A(n585), .B(n584), .ZN(n626) );
  AND2_X1 U447 ( .A1(n583), .A2(n409), .ZN(n408) );
  XNOR2_X1 U448 ( .A(n523), .B(n522), .ZN(n548) );
  XNOR2_X1 U449 ( .A(KEYINPUT13), .B(G475), .ZN(n522) );
  INV_X1 U450 ( .A(KEYINPUT19), .ZN(n414) );
  XNOR2_X1 U451 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U452 ( .A(n646), .B(KEYINPUT88), .ZN(n742) );
  INV_X1 U453 ( .A(KEYINPUT42), .ZN(n598) );
  OR2_X1 U454 ( .A1(n626), .A2(n671), .ZN(n686) );
  XOR2_X1 U455 ( .A(G131), .B(KEYINPUT4), .Z(n351) );
  XOR2_X1 U456 ( .A(n612), .B(KEYINPUT78), .Z(n352) );
  XOR2_X1 U457 ( .A(n536), .B(KEYINPUT79), .Z(n353) );
  OR2_X1 U458 ( .A1(n582), .A2(n498), .ZN(n354) );
  AND2_X1 U459 ( .A1(n552), .A2(n590), .ZN(n355) );
  AND2_X1 U460 ( .A1(n601), .A2(n704), .ZN(n356) );
  INV_X1 U461 ( .A(G101), .ZN(n423) );
  AND2_X1 U462 ( .A1(n547), .A2(n590), .ZN(n357) );
  XOR2_X1 U463 ( .A(n732), .B(n731), .Z(n358) );
  XNOR2_X1 U464 ( .A(n360), .B(KEYINPUT73), .ZN(n359) );
  NAND2_X1 U465 ( .A1(n362), .A2(n361), .ZN(n360) );
  XNOR2_X1 U466 ( .A(n620), .B(KEYINPUT47), .ZN(n361) );
  INV_X1 U467 ( .A(n674), .ZN(n362) );
  NAND2_X1 U468 ( .A1(n363), .A2(n623), .ZN(n685) );
  XNOR2_X1 U469 ( .A(n606), .B(n605), .ZN(n363) );
  INV_X1 U470 ( .A(n373), .ZN(n365) );
  NAND2_X1 U471 ( .A1(n649), .A2(n369), .ZN(n368) );
  NAND2_X1 U472 ( .A1(n373), .A2(n371), .ZN(n370) );
  AND2_X1 U473 ( .A1(n372), .A2(KEYINPUT83), .ZN(n371) );
  INV_X1 U474 ( .A(n649), .ZN(n372) );
  NAND2_X1 U475 ( .A1(n518), .A2(G210), .ZN(n375) );
  AND2_X1 U476 ( .A1(n554), .A2(n356), .ZN(n602) );
  INV_X1 U477 ( .A(n554), .ZN(n379) );
  NAND2_X2 U478 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X2 U479 ( .A(n566), .B(KEYINPUT45), .ZN(n637) );
  NOR2_X1 U480 ( .A1(n676), .A2(n695), .ZN(n620) );
  XNOR2_X2 U481 ( .A(n380), .B(G146), .ZN(n473) );
  AND2_X1 U482 ( .A1(n692), .A2(n383), .ZN(n382) );
  INV_X1 U483 ( .A(n615), .ZN(n384) );
  NAND2_X1 U484 ( .A1(n615), .A2(KEYINPUT85), .ZN(n388) );
  XNOR2_X2 U485 ( .A(n604), .B(n414), .ZN(n618) );
  NAND2_X1 U486 ( .A1(n394), .A2(n389), .ZN(n557) );
  NAND2_X1 U487 ( .A1(n400), .A2(n391), .ZN(n390) );
  NAND2_X1 U488 ( .A1(n393), .A2(KEYINPUT103), .ZN(n392) );
  INV_X1 U489 ( .A(n400), .ZN(n393) );
  NAND2_X1 U490 ( .A1(n681), .A2(n396), .ZN(n395) );
  NAND2_X1 U491 ( .A1(n398), .A2(n400), .ZN(n397) );
  NOR2_X1 U492 ( .A1(n681), .A2(n399), .ZN(n398) );
  INV_X1 U493 ( .A(KEYINPUT103), .ZN(n399) );
  NAND2_X1 U494 ( .A1(n547), .A2(n355), .ZN(n400) );
  XNOR2_X2 U495 ( .A(n401), .B(KEYINPUT35), .ZN(n653) );
  NAND2_X1 U496 ( .A1(n402), .A2(n352), .ZN(n401) );
  XNOR2_X1 U497 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U498 ( .A(KEYINPUT34), .ZN(n403) );
  NAND2_X1 U499 ( .A1(n502), .A2(n544), .ZN(n404) );
  XNOR2_X2 U500 ( .A(n406), .B(G143), .ZN(n474) );
  NAND2_X1 U501 ( .A1(n408), .A2(n609), .ZN(n585) );
  INV_X1 U502 ( .A(n611), .ZN(n410) );
  INV_X1 U503 ( .A(KEYINPUT48), .ZN(n411) );
  NAND2_X1 U504 ( .A1(n413), .A2(n607), .ZN(n412) );
  NAND2_X1 U505 ( .A1(n618), .A2(n354), .ZN(n501) );
  NAND2_X1 U506 ( .A1(n416), .A2(n353), .ZN(n537) );
  XNOR2_X2 U507 ( .A(n531), .B(n417), .ZN(n416) );
  XNOR2_X1 U508 ( .A(n456), .B(n418), .ZN(n420) );
  XNOR2_X1 U509 ( .A(n733), .B(n358), .ZN(n734) );
  NAND2_X1 U510 ( .A1(n738), .A2(G469), .ZN(n733) );
  AND2_X2 U511 ( .A1(n559), .A2(n558), .ZN(n565) );
  XOR2_X1 U512 ( .A(n430), .B(n429), .Z(n422) );
  INV_X1 U513 ( .A(KEYINPUT76), .ZN(n627) );
  XNOR2_X1 U514 ( .A(n483), .B(n422), .ZN(n431) );
  XNOR2_X1 U515 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n576) );
  XNOR2_X1 U516 ( .A(n505), .B(KEYINPUT9), .ZN(n506) );
  XNOR2_X1 U517 ( .A(n599), .B(n598), .ZN(n769) );
  XNOR2_X1 U518 ( .A(G110), .B(G104), .ZN(n424) );
  XOR2_X1 U519 ( .A(KEYINPUT89), .B(G107), .Z(n425) );
  INV_X1 U520 ( .A(KEYINPUT70), .ZN(n427) );
  XNOR2_X1 U521 ( .A(n427), .B(KEYINPUT71), .ZN(n428) );
  XOR2_X1 U522 ( .A(G146), .B(KEYINPUT93), .Z(n430) );
  NAND2_X1 U523 ( .A1(G227), .A2(n440), .ZN(n429) );
  XOR2_X1 U524 ( .A(G137), .B(G140), .Z(n442) );
  NOR2_X1 U525 ( .A1(n730), .A2(G902), .ZN(n432) );
  XNOR2_X2 U526 ( .A(n432), .B(G469), .ZN(n594) );
  INV_X1 U527 ( .A(KEYINPUT65), .ZN(n433) );
  XNOR2_X1 U528 ( .A(n433), .B(KEYINPUT1), .ZN(n434) );
  XNOR2_X1 U529 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n435) );
  XOR2_X2 U530 ( .A(n473), .B(KEYINPUT10), .Z(n760) );
  XNOR2_X1 U531 ( .A(n435), .B(n760), .ZN(n439) );
  XOR2_X1 U532 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n437) );
  XNOR2_X1 U533 ( .A(G110), .B(KEYINPUT94), .ZN(n436) );
  XNOR2_X1 U534 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U535 ( .A(n439), .B(n438), .ZN(n447) );
  NAND2_X1 U536 ( .A1(n440), .A2(G234), .ZN(n441) );
  XOR2_X1 U537 ( .A(n441), .B(KEYINPUT8), .Z(n504) );
  AND2_X1 U538 ( .A1(G221), .A2(n504), .ZN(n445) );
  XNOR2_X1 U539 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U540 ( .A(n447), .B(n446), .ZN(n739) );
  NOR2_X1 U541 ( .A1(G902), .A2(n739), .ZN(n452) );
  XOR2_X1 U542 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n450) );
  XNOR2_X1 U543 ( .A(KEYINPUT15), .B(G902), .ZN(n569) );
  NAND2_X1 U544 ( .A1(n569), .A2(G234), .ZN(n448) );
  XNOR2_X1 U545 ( .A(n448), .B(KEYINPUT20), .ZN(n453) );
  NAND2_X1 U546 ( .A1(G217), .A2(n453), .ZN(n449) );
  XNOR2_X1 U547 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X2 U548 ( .A(n452), .B(n451), .ZN(n703) );
  NAND2_X1 U549 ( .A1(n453), .A2(G221), .ZN(n455) );
  INV_X1 U550 ( .A(KEYINPUT21), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n455), .B(n454), .ZN(n704) );
  NAND2_X1 U552 ( .A1(n703), .A2(n704), .ZN(n700) );
  XNOR2_X1 U553 ( .A(KEYINPUT90), .B(KEYINPUT3), .ZN(n456) );
  INV_X1 U554 ( .A(KEYINPUT5), .ZN(n457) );
  INV_X1 U555 ( .A(n464), .ZN(n462) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT75), .Z(n459) );
  XNOR2_X1 U557 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U558 ( .A(n460), .B(G137), .ZN(n463) );
  INV_X1 U559 ( .A(n463), .ZN(n461) );
  NAND2_X1 U560 ( .A1(n462), .A2(n461), .ZN(n466) );
  NAND2_X1 U561 ( .A1(n464), .A2(n463), .ZN(n465) );
  INV_X1 U562 ( .A(G902), .ZN(n486) );
  XNOR2_X1 U563 ( .A(KEYINPUT101), .B(G472), .ZN(n468) );
  XNOR2_X2 U564 ( .A(n469), .B(n468), .ZN(n590) );
  XNOR2_X1 U565 ( .A(n590), .B(KEYINPUT6), .ZN(n554) );
  INV_X1 U566 ( .A(n720), .ZN(n502) );
  XNOR2_X1 U567 ( .A(KEYINPUT16), .B(G122), .ZN(n470) );
  XNOR2_X1 U568 ( .A(n470), .B(KEYINPUT72), .ZN(n471) );
  XNOR2_X1 U569 ( .A(KEYINPUT4), .B(n473), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U571 ( .A(n477), .B(n476), .ZN(n481) );
  NAND2_X1 U572 ( .A1(G224), .A2(n440), .ZN(n479) );
  XOR2_X1 U573 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n478) );
  XNOR2_X1 U574 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U575 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U576 ( .A(n751), .B(n482), .ZN(n484) );
  XNOR2_X1 U577 ( .A(n484), .B(n483), .ZN(n640) );
  NAND2_X1 U578 ( .A1(n640), .A2(n569), .ZN(n490) );
  NAND2_X1 U579 ( .A1(n486), .A2(n485), .ZN(n491) );
  NAND2_X1 U580 ( .A1(n491), .A2(G210), .ZN(n488) );
  INV_X1 U581 ( .A(KEYINPUT91), .ZN(n487) );
  XNOR2_X1 U582 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X2 U583 ( .A(n490), .B(n489), .ZN(n615) );
  NAND2_X1 U584 ( .A1(n491), .A2(G214), .ZN(n692) );
  XNOR2_X1 U585 ( .A(n492), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U586 ( .A1(n493), .A2(G952), .ZN(n719) );
  NOR2_X1 U587 ( .A1(n719), .A2(G953), .ZN(n582) );
  NAND2_X1 U588 ( .A1(n493), .A2(G902), .ZN(n577) );
  INV_X1 U589 ( .A(n577), .ZN(n495) );
  INV_X1 U590 ( .A(G953), .ZN(n494) );
  NOR2_X1 U591 ( .A1(G898), .A2(n494), .ZN(n753) );
  NAND2_X1 U592 ( .A1(n495), .A2(n753), .ZN(n497) );
  INV_X1 U593 ( .A(KEYINPUT92), .ZN(n496) );
  XNOR2_X1 U594 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U595 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n499) );
  XNOR2_X1 U596 ( .A(n499), .B(KEYINPUT67), .ZN(n500) );
  XNOR2_X2 U597 ( .A(n501), .B(n500), .ZN(n544) );
  INV_X1 U598 ( .A(n503), .ZN(n511) );
  NAND2_X1 U599 ( .A1(G217), .A2(n504), .ZN(n507) );
  XOR2_X1 U600 ( .A(G107), .B(KEYINPUT7), .Z(n505) );
  XOR2_X1 U601 ( .A(G116), .B(G122), .Z(n508) );
  XNOR2_X1 U602 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n511), .B(n510), .ZN(n735) );
  XOR2_X1 U604 ( .A(G478), .B(n529), .Z(n551) );
  XNOR2_X1 U605 ( .A(G113), .B(G131), .ZN(n512) );
  XNOR2_X1 U606 ( .A(n513), .B(n512), .ZN(n517) );
  XOR2_X1 U607 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n515) );
  XNOR2_X1 U608 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U609 ( .A(n517), .B(n516), .Z(n521) );
  NAND2_X1 U610 ( .A1(G214), .A2(n518), .ZN(n519) );
  XNOR2_X1 U611 ( .A(n760), .B(n519), .ZN(n520) );
  XNOR2_X1 U612 ( .A(n521), .B(n520), .ZN(n656) );
  NOR2_X1 U613 ( .A1(G902), .A2(n656), .ZN(n523) );
  NAND2_X1 U614 ( .A1(n551), .A2(n548), .ZN(n612) );
  INV_X1 U615 ( .A(n653), .ZN(n560) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n524) );
  AND2_X1 U617 ( .A1(n524), .A2(KEYINPUT68), .ZN(n525) );
  NAND2_X1 U618 ( .A1(n560), .A2(n525), .ZN(n528) );
  INV_X1 U619 ( .A(KEYINPUT68), .ZN(n526) );
  NAND2_X1 U620 ( .A1(n653), .A2(n526), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n528), .A2(n527), .ZN(n538) );
  XNOR2_X1 U622 ( .A(G478), .B(n529), .ZN(n549) );
  INV_X1 U623 ( .A(n548), .ZN(n550) );
  NAND2_X1 U624 ( .A1(n549), .A2(n550), .ZN(n587) );
  INV_X1 U625 ( .A(n704), .ZN(n589) );
  NOR2_X1 U626 ( .A1(n587), .A2(n589), .ZN(n530) );
  NAND2_X1 U627 ( .A1(n544), .A2(n530), .ZN(n531) );
  INV_X1 U628 ( .A(n701), .ZN(n623) );
  INV_X1 U629 ( .A(n703), .ZN(n574) );
  AND2_X1 U630 ( .A1(n590), .A2(n574), .ZN(n532) );
  NOR2_X1 U631 ( .A1(n701), .A2(n703), .ZN(n534) );
  XOR2_X1 U632 ( .A(KEYINPUT104), .B(n534), .Z(n535) );
  NOR2_X1 U633 ( .A1(n535), .A2(n554), .ZN(n536) );
  XNOR2_X1 U634 ( .A(n537), .B(KEYINPUT32), .ZN(n652) );
  NAND2_X1 U635 ( .A1(n561), .A2(n538), .ZN(n559) );
  INV_X1 U636 ( .A(n539), .ZN(n540) );
  INV_X1 U637 ( .A(n590), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n540), .A2(n575), .ZN(n541) );
  XNOR2_X1 U639 ( .A(n541), .B(KEYINPUT102), .ZN(n709) );
  INV_X1 U640 ( .A(n709), .ZN(n542) );
  NAND2_X1 U641 ( .A1(n542), .A2(n544), .ZN(n543) );
  NOR2_X1 U642 ( .A1(n594), .A2(n700), .ZN(n608) );
  NAND2_X1 U643 ( .A1(n544), .A2(n608), .ZN(n546) );
  INV_X1 U644 ( .A(KEYINPUT98), .ZN(n545) );
  XNOR2_X1 U645 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U646 ( .A1(n549), .A2(n548), .ZN(n675) );
  NAND2_X1 U647 ( .A1(n551), .A2(n550), .ZN(n671) );
  AND2_X1 U648 ( .A1(n675), .A2(n671), .ZN(n695) );
  INV_X1 U649 ( .A(n695), .ZN(n552) );
  INV_X1 U650 ( .A(n553), .ZN(n556) );
  NOR2_X1 U651 ( .A1(n554), .A2(n574), .ZN(n555) );
  AND2_X1 U652 ( .A1(n556), .A2(n555), .ZN(n651) );
  NOR2_X1 U653 ( .A1(n557), .A2(n651), .ZN(n558) );
  AND2_X1 U654 ( .A1(n560), .A2(KEYINPUT68), .ZN(n562) );
  NAND2_X1 U655 ( .A1(n561), .A2(n562), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n563), .A2(KEYINPUT44), .ZN(n564) );
  INV_X1 U657 ( .A(KEYINPUT2), .ZN(n567) );
  NOR2_X1 U658 ( .A1(n567), .A2(KEYINPUT82), .ZN(n568) );
  NAND2_X1 U659 ( .A1(n569), .A2(n568), .ZN(n631) );
  INV_X1 U660 ( .A(n631), .ZN(n571) );
  INV_X1 U661 ( .A(n569), .ZN(n570) );
  OR2_X1 U662 ( .A1(n571), .A2(n570), .ZN(n630) );
  AND2_X1 U663 ( .A1(n637), .A2(n630), .ZN(n629) );
  INV_X1 U664 ( .A(n594), .ZN(n572) );
  NAND2_X1 U665 ( .A1(n704), .A2(n572), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n583) );
  XNOR2_X1 U667 ( .A(n615), .B(KEYINPUT38), .ZN(n691) );
  NOR2_X1 U668 ( .A1(n440), .A2(n577), .ZN(n578) );
  XOR2_X1 U669 ( .A(KEYINPUT106), .B(n578), .Z(n579) );
  NOR2_X1 U670 ( .A1(G900), .A2(n579), .ZN(n580) );
  XOR2_X1 U671 ( .A(KEYINPUT107), .B(n580), .Z(n581) );
  NOR2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n611) );
  XOR2_X1 U673 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n584) );
  XNOR2_X1 U674 ( .A(n586), .B(KEYINPUT40), .ZN(n770) );
  NAND2_X1 U675 ( .A1(n691), .A2(n692), .ZN(n694) );
  INV_X1 U676 ( .A(n721), .ZN(n597) );
  NOR2_X1 U677 ( .A1(n703), .A2(n611), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n590), .A2(n589), .ZN(n591) );
  AND2_X1 U679 ( .A1(n601), .A2(n591), .ZN(n593) );
  XNOR2_X1 U680 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n592) );
  XNOR2_X1 U681 ( .A(n593), .B(n592), .ZN(n596) );
  XNOR2_X1 U682 ( .A(KEYINPUT110), .B(n594), .ZN(n595) );
  NAND2_X1 U683 ( .A1(n597), .A2(n619), .ZN(n599) );
  NOR2_X1 U684 ( .A1(n770), .A2(n769), .ZN(n600) );
  XNOR2_X1 U685 ( .A(n600), .B(KEYINPUT46), .ZN(n607) );
  XOR2_X1 U686 ( .A(KEYINPUT108), .B(n602), .Z(n603) );
  NOR2_X1 U687 ( .A1(n603), .A2(n675), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n621), .A2(n604), .ZN(n606) );
  XOR2_X1 U689 ( .A(KEYINPUT36), .B(KEYINPUT112), .Z(n605) );
  NAND2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n614) );
  INV_X1 U692 ( .A(n612), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n617) );
  BUF_X1 U694 ( .A(n615), .Z(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n674) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n676) );
  NAND2_X1 U697 ( .A1(n621), .A2(n692), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT43), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n625), .A2(n384), .ZN(n649) );
  XNOR2_X1 U701 ( .A(n765), .B(n627), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n636) );
  INV_X1 U703 ( .A(n630), .ZN(n634) );
  NAND2_X1 U704 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n632) );
  AND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  OR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n639) );
  INV_X1 U708 ( .A(n637), .ZN(n743) );
  NOR2_X2 U709 ( .A1(n743), .A2(n765), .ZN(n690) );
  NAND2_X1 U710 ( .A1(n690), .A2(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n729), .A2(G210), .ZN(n645) );
  XOR2_X1 U712 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n642) );
  XNOR2_X1 U713 ( .A(KEYINPUT80), .B(KEYINPUT55), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n640), .B(n643), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n647) );
  NOR2_X1 U717 ( .A1(n440), .A2(G952), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n648), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U719 ( .A(G140), .B(n649), .Z(G42) );
  INV_X1 U720 ( .A(n675), .ZN(n678) );
  NAND2_X1 U721 ( .A1(n357), .A2(n678), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n650), .B(n347), .ZN(G6) );
  XOR2_X1 U723 ( .A(G101), .B(n651), .Z(G3) );
  XNOR2_X1 U724 ( .A(n652), .B(G119), .ZN(G21) );
  XOR2_X1 U725 ( .A(G122), .B(n653), .Z(G24) );
  XNOR2_X1 U726 ( .A(G110), .B(KEYINPUT114), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n350), .B(n654), .ZN(G12) );
  NAND2_X1 U728 ( .A1(n729), .A2(G475), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT59), .B(n656), .Z(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(G60) );
  XOR2_X1 U733 ( .A(n662), .B(KEYINPUT62), .Z(n663) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT63), .B(KEYINPUT113), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(G57) );
  INV_X1 U737 ( .A(n671), .ZN(n680) );
  NAND2_X1 U738 ( .A1(n357), .A2(n680), .ZN(n669) );
  XOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U741 ( .A(G107), .B(n670), .ZN(G9) );
  NOR2_X1 U742 ( .A1(n676), .A2(n671), .ZN(n673) );
  XNOR2_X1 U743 ( .A(G128), .B(KEYINPUT29), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(G30) );
  XOR2_X1 U745 ( .A(G143), .B(n674), .Z(G45) );
  NOR2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U747 ( .A(G146), .B(n677), .Z(G48) );
  NAND2_X1 U748 ( .A1(n681), .A2(n678), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(G113), .ZN(G15) );
  XOR2_X1 U750 ( .A(G116), .B(KEYINPUT115), .Z(n683) );
  NAND2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(G18) );
  XOR2_X1 U753 ( .A(G125), .B(KEYINPUT37), .Z(n684) );
  XNOR2_X1 U754 ( .A(n685), .B(n684), .ZN(G27) );
  INV_X1 U755 ( .A(n686), .ZN(n687) );
  XOR2_X1 U756 ( .A(G134), .B(n687), .Z(n688) );
  XNOR2_X1 U757 ( .A(KEYINPUT116), .B(n688), .ZN(G36) );
  XOR2_X1 U758 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n689) );
  XNOR2_X1 U759 ( .A(n690), .B(n689), .ZN(n725) );
  NOR2_X1 U760 ( .A1(n691), .A2(n692), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n587), .A2(n693), .ZN(n697) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U764 ( .A1(n720), .A2(n698), .ZN(n715) );
  XNOR2_X1 U765 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT51), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U768 ( .A(KEYINPUT50), .B(n702), .ZN(n708) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U770 ( .A(KEYINPUT49), .B(n705), .Z(n706) );
  NOR2_X1 U771 ( .A1(n575), .A2(n706), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U774 ( .A(n712), .B(n711), .Z(n713) );
  NOR2_X1 U775 ( .A1(n721), .A2(n713), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U777 ( .A(KEYINPUT52), .B(n716), .Z(n717) );
  XNOR2_X1 U778 ( .A(n717), .B(KEYINPUT119), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U781 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U782 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U783 ( .A(KEYINPUT120), .B(n726), .ZN(n727) );
  NOR2_X2 U784 ( .A1(n727), .A2(G953), .ZN(n728) );
  XNOR2_X1 U785 ( .A(n728), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U786 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n732) );
  XNOR2_X1 U787 ( .A(n730), .B(KEYINPUT57), .ZN(n731) );
  NOR2_X1 U788 ( .A1(n742), .A2(n734), .ZN(G54) );
  NAND2_X1 U789 ( .A1(n738), .A2(G478), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U791 ( .A1(n742), .A2(n737), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n738), .A2(G217), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U794 ( .A1(n742), .A2(n741), .ZN(G66) );
  NOR2_X1 U795 ( .A1(n743), .A2(G953), .ZN(n750) );
  XOR2_X1 U796 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n745) );
  NAND2_X1 U797 ( .A1(G224), .A2(G953), .ZN(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U799 ( .A(KEYINPUT123), .B(n746), .ZN(n747) );
  NAND2_X1 U800 ( .A1(n747), .A2(G898), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(KEYINPUT125), .ZN(n749) );
  NOR2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n758) );
  XNOR2_X1 U803 ( .A(n752), .B(n751), .ZN(n755) );
  INV_X1 U804 ( .A(n753), .ZN(n754) );
  AND2_X1 U805 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U806 ( .A(KEYINPUT126), .B(n756), .Z(n757) );
  XNOR2_X1 U807 ( .A(n758), .B(n757), .ZN(G69) );
  XOR2_X1 U808 ( .A(n760), .B(n759), .Z(n764) );
  XOR2_X1 U809 ( .A(G227), .B(n764), .Z(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n762), .A2(G953), .ZN(n763) );
  XOR2_X1 U812 ( .A(KEYINPUT127), .B(n763), .Z(n768) );
  XOR2_X1 U813 ( .A(n765), .B(n764), .Z(n766) );
  NAND2_X1 U814 ( .A1(n766), .A2(n440), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n768), .A2(n767), .ZN(G72) );
  XOR2_X1 U816 ( .A(n769), .B(G137), .Z(G39) );
  XOR2_X1 U817 ( .A(G131), .B(n770), .Z(G33) );
endmodule

