//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n206), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n214), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT67), .Z(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  AND2_X1   g0034(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n225), .A2(new_n234), .A3(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n220), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n208), .A2(G20), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  NAND2_X1  g0057(.A1(new_n212), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n255), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n211), .A2(KEYINPUT69), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G1), .ZN(new_n266));
  AOI211_X1 g0066(.A(new_n263), .B(new_n212), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n212), .B1(new_n264), .B2(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n266), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n255), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(KEYINPUT71), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n255), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT72), .B(new_n269), .C1(new_n277), .C2(new_n207), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n207), .B1(new_n274), .B2(new_n276), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n268), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n262), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n211), .B(G274), .C1(G41), .C2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n289), .B1(new_n290), .B2(new_n287), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n220), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n286), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G41), .A2(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n264), .B2(new_n266), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT70), .B1(new_n298), .B2(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  INV_X1    g0100(.A(G33), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  OAI211_X1 g0102(.A(G1), .B(G13), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT69), .B(G1), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n303), .C1(new_n304), .C2(new_n297), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G226), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(KEYINPUT73), .B(G200), .Z(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n308), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n282), .B2(KEYINPUT9), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT10), .B1(new_n284), .B2(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n283), .A4(new_n312), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n278), .A2(new_n281), .ZN(new_n319));
  INV_X1    g0119(.A(new_n262), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n308), .A2(G179), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n308), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT75), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n299), .A2(G238), .A3(new_n305), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT74), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(G33), .A3(G97), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G33), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n335), .A3(G232), .A4(G1698), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(G226), .A4(new_n288), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n295), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n327), .A2(new_n339), .A3(new_n285), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT13), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n327), .A2(new_n339), .A3(new_n342), .A4(new_n285), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(G190), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n272), .A2(G68), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n260), .A2(G50), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n347), .B1(new_n212), .B2(G68), .C1(new_n290), .C2(new_n258), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n254), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n270), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G68), .A3(new_n255), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n344), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n341), .B2(new_n343), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n326), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n341), .A2(new_n343), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G200), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n356), .A4(new_n344), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n356), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(G169), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n361), .A2(new_n368), .A3(G169), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n341), .A2(G179), .A3(new_n343), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n364), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT71), .B1(new_n267), .B2(new_n254), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(new_n257), .A3(new_n352), .A4(new_n276), .ZN(new_n375));
  INV_X1    g0175(.A(new_n257), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n267), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n287), .B2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n333), .A2(new_n335), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n202), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n203), .A2(new_n205), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n260), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n379), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(new_n254), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n382), .B2(new_n212), .ZN(new_n392));
  AOI211_X1 g0192(.A(new_n380), .B(G20), .C1(new_n333), .C2(new_n335), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n378), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n333), .A2(new_n335), .A3(G223), .A4(new_n288), .ZN(new_n398));
  INV_X1    g0198(.A(G87), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n301), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n287), .A2(G226), .A3(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n295), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(G232), .B(new_n303), .C1(new_n304), .C2(new_n297), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT76), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n286), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n298), .A2(new_n295), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT76), .A3(G232), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n323), .ZN(new_n409));
  INV_X1    g0209(.A(G179), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n402), .A2(new_n405), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n373), .B1(new_n397), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n409), .A2(new_n411), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n375), .A2(new_n377), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n396), .A2(new_n390), .A3(new_n254), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(G200), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n402), .A2(new_n405), .A3(new_n407), .A4(G190), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n397), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n415), .A2(new_n416), .A3(new_n419), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n413), .A2(new_n418), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n306), .A2(G244), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n428));
  INV_X1    g0228(.A(G107), .ZN(new_n429));
  INV_X1    g0229(.A(G238), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n428), .B1(new_n429), .B2(new_n287), .C1(new_n291), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n295), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n285), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n311), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n352), .A2(G77), .A3(new_n255), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G77), .B2(new_n272), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n257), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n437));
  XOR2_X1   g0237(.A(KEYINPUT15), .B(G87), .Z(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n259), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n255), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n434), .B(new_n441), .C1(new_n309), .C2(new_n433), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n433), .B2(new_n323), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G179), .B2(new_n433), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n426), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AND4_X1   g0245(.A1(new_n318), .A2(new_n325), .A3(new_n372), .A4(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n333), .A2(new_n335), .A3(G264), .A4(G1698), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT81), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n287), .A2(KEYINPUT81), .A3(G264), .A4(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n382), .A2(G303), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n287), .A2(G257), .A3(new_n288), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n295), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n264), .B2(new_n266), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n295), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G274), .B1(new_n294), .B2(new_n220), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n459), .A2(new_n304), .A3(new_n455), .ZN(new_n460));
  AOI22_X1  g0260(.A1(G270), .A2(new_n458), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G169), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n212), .C1(G33), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G20), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT82), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n253), .A2(new_n220), .B1(G20), .B2(new_n468), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n467), .A4(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT83), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n467), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(KEYINPUT83), .B(KEYINPUT20), .C1(new_n472), .C2(new_n467), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n475), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n272), .A2(G116), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n271), .A2(G33), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n272), .A2(new_n255), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n468), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n464), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n477), .A2(new_n478), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT83), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n477), .A2(new_n476), .A3(new_n478), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n474), .A3(new_n471), .A4(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n272), .A2(new_n255), .A3(new_n484), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n482), .B1(new_n492), .B2(G116), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT84), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n463), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT84), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT84), .B1(new_n491), .B2(new_n493), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n323), .B1(new_n454), .B2(new_n461), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n271), .A2(G45), .ZN(new_n502));
  INV_X1    g0302(.A(new_n457), .ZN(new_n503));
  OAI211_X1 g0303(.A(G270), .B(new_n303), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n456), .A2(G274), .A3(new_n303), .A4(new_n457), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n295), .B2(new_n453), .ZN(new_n507));
  AOI22_X1  g0307(.A1(KEYINPUT21), .A2(new_n501), .B1(new_n507), .B2(G179), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n495), .A2(new_n497), .B1(new_n500), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n462), .A2(G200), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n309), .B2(new_n462), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n499), .A3(new_n498), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n333), .A2(new_n335), .A3(G250), .A4(new_n288), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT86), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n287), .A2(KEYINPUT86), .A3(G250), .A4(new_n288), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G294), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n287), .A2(G257), .A3(G1698), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n295), .ZN(new_n521));
  AOI22_X1  g0321(.A1(G264), .A2(new_n458), .B1(new_n460), .B2(new_n457), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n410), .ZN(new_n523));
  OAI211_X1 g0323(.A(G264), .B(new_n303), .C1(new_n502), .C2(new_n503), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n505), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n295), .B2(new_n520), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n526), .B2(G169), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n492), .A2(G107), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n272), .B2(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n429), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n333), .A2(new_n335), .A3(new_n212), .A4(G87), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n287), .A2(new_n536), .A3(new_n212), .A4(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G116), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n212), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n429), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT24), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n255), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n544), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n535), .B2(new_n537), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n533), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n527), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n521), .A2(new_n522), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n521), .A2(new_n522), .A3(G190), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(G107), .A2(new_n492), .B1(new_n530), .B2(new_n531), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n254), .B1(new_n549), .B2(KEYINPUT24), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n545), .A2(new_n546), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n553), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n551), .A2(KEYINPUT87), .A3(new_n556), .A4(new_n555), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n552), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n267), .A2(new_n466), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n492), .A2(G97), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n429), .B1(new_n381), .B2(new_n383), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n466), .A2(new_n429), .A3(KEYINPUT6), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n429), .A2(KEYINPUT77), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G107), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n568), .A2(new_n570), .A3(new_n572), .A4(new_n574), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n212), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n260), .A2(G77), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n567), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n565), .B(new_n566), .C1(new_n581), .C2(new_n255), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n333), .A2(new_n335), .A3(G244), .A4(new_n288), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n465), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n295), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n458), .A2(G257), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n505), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n323), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n588), .A2(new_n295), .B1(G257), .B2(new_n458), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n410), .A3(new_n505), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n582), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n271), .A2(new_n303), .A3(G45), .A4(G274), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n303), .B1(new_n304), .B2(new_n455), .ZN(new_n597));
  INV_X1    g0397(.A(G250), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n333), .A2(new_n335), .A3(G238), .A4(new_n288), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT78), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n287), .A2(new_n602), .A3(G238), .A4(new_n288), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n287), .A2(G244), .A3(G1698), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n601), .A2(new_n603), .A3(new_n539), .A4(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(G179), .B(new_n599), .C1(new_n295), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n295), .ZN(new_n607));
  INV_X1    g0407(.A(new_n599), .ZN(new_n608));
  AOI21_X1  g0408(.A(G169), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  INV_X1    g0411(.A(new_n438), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n485), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n254), .B1(new_n270), .B2(G13), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(KEYINPUT79), .A3(new_n438), .A4(new_n484), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n399), .A2(new_n466), .A3(new_n429), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n329), .B2(new_n331), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(G20), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n333), .A2(new_n335), .A3(new_n212), .A4(G68), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n258), .B2(new_n466), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n255), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n272), .A2(new_n438), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT80), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n616), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n616), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n610), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n591), .A2(G200), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n565), .B1(new_n485), .B2(new_n466), .ZN(new_n632));
  INV_X1    g0432(.A(new_n578), .ZN(new_n633));
  OAI21_X1  g0433(.A(G107), .B1(new_n392), .B2(new_n393), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(new_n579), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n254), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n593), .A2(G190), .A3(new_n505), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n485), .A2(new_n399), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n624), .A2(new_n639), .A3(new_n625), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n599), .B1(new_n605), .B2(new_n295), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G190), .ZN(new_n642));
  INV_X1    g0442(.A(new_n311), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n642), .C1(new_n643), .C2(new_n641), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n595), .A2(new_n630), .A3(new_n638), .A4(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n446), .A2(new_n513), .A3(new_n564), .A4(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n325), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n423), .A2(new_n425), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n371), .A2(new_n365), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n362), .A2(new_n356), .A3(new_n344), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n650), .B(new_n443), .C1(G179), .C2(new_n433), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n413), .A2(new_n418), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(KEYINPUT90), .B1(new_n314), .B2(new_n317), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT90), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n652), .B2(new_n653), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n562), .A2(new_n563), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n595), .A2(new_n638), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n626), .B1(new_n399), .B2(new_n485), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n641), .A2(new_n643), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT88), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n640), .B(new_n664), .C1(new_n643), .C2(new_n641), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n665), .A3(new_n642), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n659), .A2(new_n660), .A3(new_n630), .A4(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT89), .B1(new_n527), .B2(new_n551), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n554), .A2(new_n323), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n561), .A2(new_n669), .A3(new_n670), .A4(new_n523), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n509), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n582), .A2(new_n592), .A3(new_n594), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n630), .A2(new_n675), .A3(new_n644), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n666), .A2(new_n678), .A3(new_n675), .A4(new_n630), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n679), .A3(new_n630), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n446), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n658), .A2(new_n681), .ZN(G369));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  XNOR2_X1  g0483(.A(KEYINPUT91), .B(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n212), .A2(G13), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n304), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n304), .B2(new_n685), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT92), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n686), .A2(new_n690), .A3(G213), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n513), .B1(new_n500), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n509), .B(new_n694), .C1(new_n499), .C2(new_n498), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n683), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n564), .B1(new_n551), .B2(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n509), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n552), .A2(new_n694), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n564), .A2(new_n509), .A3(new_n695), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n672), .A2(new_n695), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n215), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n617), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n219), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n711), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n593), .A2(new_n521), .A3(new_n522), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n454), .A2(new_n461), .A3(G179), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n641), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n593), .A2(new_n641), .A3(new_n521), .A4(new_n522), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n718), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n607), .A2(new_n608), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n641), .A2(KEYINPUT93), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n591), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n462), .A2(new_n554), .A3(new_n410), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n694), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT31), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n734), .B(new_n694), .C1(new_n724), .C2(new_n731), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n513), .A2(new_n645), .A3(new_n564), .A4(new_n695), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n683), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n667), .A2(new_n673), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n677), .A2(new_n630), .A3(new_n679), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n694), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n630), .A2(new_n675), .A3(new_n678), .A4(new_n644), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(new_n630), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n666), .A2(new_n675), .A3(new_n630), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT26), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n509), .A2(new_n552), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n744), .B(new_n746), .C1(new_n667), .C2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n738), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n716), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(new_n698), .ZN(new_n752));
  INV_X1    g0552(.A(new_n685), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n211), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n710), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n696), .A2(new_n683), .A3(new_n697), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n752), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n696), .A2(new_n697), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n215), .A2(new_n287), .ZN(new_n764));
  INV_X1    g0564(.A(G355), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n765), .B1(G116), .B2(new_n215), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n248), .A2(G45), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n709), .A2(new_n287), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n219), .B2(new_n455), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n220), .B1(G20), .B2(new_n323), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n756), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n410), .A2(new_n358), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n212), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n212), .A2(new_n309), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n410), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G322), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n778), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G179), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n778), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n780), .B(new_n787), .C1(G329), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n781), .A2(new_n777), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT95), .B(G326), .Z(new_n794));
  AOI21_X1  g0594(.A(new_n212), .B1(new_n788), .B2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n793), .A2(new_n794), .B1(new_n796), .B2(G294), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n311), .A2(new_n410), .A3(new_n778), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G283), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n791), .A2(new_n798), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n311), .A2(new_n410), .A3(new_n781), .ZN(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n382), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n792), .A2(new_n207), .B1(new_n779), .B2(new_n202), .ZN(new_n808));
  INV_X1    g0608(.A(new_n785), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G77), .B2(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n399), .B2(new_n804), .C1(new_n429), .C2(new_n800), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n789), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n783), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n382), .B1(new_n816), .B2(G58), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(new_n466), .C2(new_n795), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n803), .A2(new_n807), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n775), .B1(new_n772), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n763), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n759), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NOR2_X1   g0623(.A1(new_n444), .A2(new_n694), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n442), .B1(new_n441), .B2(new_n695), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n444), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n741), .B(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n738), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n756), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n772), .A2(new_n760), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n757), .B1(new_n290), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n772), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n399), .A2(new_n800), .B1(new_n804), .B2(new_n429), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n382), .B1(new_n795), .B2(new_n466), .C1(new_n792), .C2(new_n805), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n785), .A2(new_n468), .B1(new_n789), .B2(new_n786), .ZN(new_n836));
  INV_X1    g0636(.A(G283), .ZN(new_n837));
  INV_X1    g0637(.A(G294), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n837), .A2(new_n779), .B1(new_n783), .B2(new_n838), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n779), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G143), .A2(new_n816), .B1(new_n841), .B2(G150), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n792), .C1(new_n812), .C2(new_n785), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n287), .B1(new_n795), .B2(new_n201), .C1(new_n846), .C2(new_n789), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n800), .A2(new_n202), .ZN(new_n848));
  INV_X1    g0648(.A(new_n804), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n847), .B(new_n848), .C1(G50), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n840), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n832), .B1(new_n833), .B2(new_n851), .C1(new_n826), .C2(new_n761), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n830), .A2(new_n852), .ZN(G384));
  NAND2_X1  g0653(.A1(new_n576), .A2(new_n577), .ZN(new_n854));
  OAI211_X1 g0654(.A(G116), .B(new_n221), .C1(new_n854), .C2(KEYINPUT35), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(KEYINPUT35), .B2(new_n854), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n219), .A2(G77), .A3(new_n385), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n207), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(G13), .B(new_n271), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT40), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n692), .B1(new_n415), .B2(new_n416), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(KEYINPUT37), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n414), .A2(new_n417), .ZN(new_n870));
  INV_X1    g0670(.A(new_n692), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n417), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n872), .A3(new_n424), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n867), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n426), .B2(new_n872), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n867), .B2(new_n869), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n863), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n876), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n864), .B1(new_n653), .B2(new_n648), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT38), .A4(new_n874), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n825), .A2(new_n444), .ZN(new_n882));
  INV_X1    g0682(.A(new_n824), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n736), .B2(new_n737), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n365), .B(new_n694), .C1(new_n364), .C2(new_n371), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n365), .A2(new_n694), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n650), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n649), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT98), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n886), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n862), .B1(new_n881), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n736), .A2(new_n737), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n870), .A2(new_n872), .A3(new_n896), .A4(new_n424), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n897), .A2(new_n898), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n879), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n863), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n880), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n886), .A2(new_n889), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT98), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT40), .A4(new_n885), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n894), .A2(new_n446), .A3(new_n895), .A4(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n894), .A2(G330), .A3(new_n910), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n446), .A2(new_n738), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n446), .B(new_n749), .C1(KEYINPUT29), .C2(new_n741), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n658), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n916), .B(new_n918), .Z(new_n919));
  OAI211_X1 g0719(.A(new_n695), .B(new_n826), .C1(new_n674), .C2(new_n680), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n883), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n877), .A2(new_n880), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(new_n909), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n653), .A2(new_n692), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n371), .A2(new_n365), .A3(new_n695), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT101), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT103), .B1(new_n903), .B2(new_n863), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT39), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n904), .A2(new_n880), .A3(KEYINPUT103), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n919), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n271), .B2(new_n753), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n919), .A2(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n861), .B1(new_n936), .B2(new_n937), .ZN(G367));
  NAND2_X1  g0738(.A1(new_n694), .A2(new_n582), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n660), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n675), .A2(new_n694), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n703), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT104), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n942), .A2(new_n509), .A3(new_n564), .A4(new_n695), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n660), .A2(new_n552), .A3(new_n939), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n694), .B1(new_n949), .B2(new_n595), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n946), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g0752(.A(KEYINPUT104), .B(new_n950), .C1(new_n947), .C2(KEYINPUT42), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(KEYINPUT42), .B2(new_n947), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n694), .A2(new_n661), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n666), .A2(new_n630), .A3(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n630), .A2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n954), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n954), .B2(new_n955), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT43), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n948), .A2(new_n951), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT104), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n948), .A2(new_n946), .A3(new_n951), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n959), .B1(new_n969), .B2(KEYINPUT105), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n954), .A2(new_n955), .A3(new_n960), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n945), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n974), .A3(new_n971), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n961), .A2(new_n962), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n944), .B(new_n975), .C1(new_n976), .C2(new_n964), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n742), .A2(new_n749), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n828), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n706), .A2(new_n943), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT107), .Z(new_n984));
  NAND3_X1  g0784(.A1(new_n707), .A2(new_n942), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n706), .B2(new_n943), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n982), .A2(new_n703), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n698), .A2(new_n702), .ZN(new_n989));
  INV_X1    g0789(.A(new_n704), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n698), .B2(new_n702), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n979), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n710), .B(KEYINPUT41), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n754), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n973), .A2(new_n977), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n769), .A2(new_n243), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n773), .B1(new_n215), .B2(new_n612), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n756), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n795), .A2(new_n202), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n779), .A2(new_n812), .B1(new_n785), .B2(new_n207), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT110), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n793), .A2(G143), .B1(new_n790), .B2(G137), .ZN(new_n1004));
  INV_X1    g0804(.A(G150), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n287), .C1(new_n1005), .C2(new_n783), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n201), .A2(new_n804), .B1(new_n800), .B2(new_n290), .ZN(new_n1007));
  OR4_X1    g0807(.A1(new_n1001), .A2(new_n1003), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n849), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT46), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n804), .B2(new_n468), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(new_n838), .C2(new_n779), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(KEYINPUT109), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT109), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G303), .A2(new_n816), .B1(new_n790), .B2(G317), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n837), .B2(new_n785), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n800), .A2(new_n466), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n382), .B1(new_n795), .B2(new_n429), .C1(new_n792), .C2(new_n786), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1008), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT47), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n833), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1000), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n762), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n959), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n997), .A2(new_n1027), .ZN(G387));
  NOR2_X1   g0828(.A1(new_n376), .A2(G50), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT50), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n712), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n455), .B1(new_n202), .B2(new_n290), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n768), .B1(new_n240), .B2(new_n455), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(G107), .B2(new_n215), .C1(new_n712), .C2(new_n764), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1037), .A2(new_n773), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n287), .B1(new_n790), .B2(new_n794), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT114), .B(G322), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n792), .A2(new_n1040), .B1(new_n779), .B2(new_n786), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT115), .ZN(new_n1042));
  INV_X1    g0842(.A(G317), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1042), .B1(new_n805), .B2(new_n785), .C1(new_n1043), .C2(new_n783), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT48), .Z(new_n1045));
  OAI22_X1  g0845(.A1(new_n804), .A2(new_n838), .B1(new_n837), .B2(new_n795), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1039), .B1(new_n468), .B2(new_n800), .C1(new_n1047), .C2(KEYINPUT49), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n849), .A2(G77), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1005), .B2(new_n789), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n382), .B(new_n1017), .C1(new_n1051), .C2(KEYINPUT112), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(KEYINPUT112), .B2(new_n1051), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT113), .Z(new_n1054));
  AOI22_X1  g0854(.A1(G50), .A2(new_n816), .B1(new_n841), .B2(new_n257), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n793), .A2(G159), .B1(new_n809), .B2(G68), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n612), .C2(new_n795), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1048), .A2(new_n1049), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n757), .B(new_n1038), .C1(new_n1058), .C2(new_n772), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n699), .A2(new_n701), .A3(new_n762), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n755), .B2(new_n992), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n710), .B(KEYINPUT116), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n750), .B2(new_n992), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT117), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n992), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n979), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1063), .B2(KEYINPUT117), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1061), .B1(new_n1064), .B2(new_n1067), .ZN(G393));
  AND3_X1   g0868(.A1(new_n978), .A2(new_n992), .A3(new_n828), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n988), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1062), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n703), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n980), .B(KEYINPUT44), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n985), .A2(new_n987), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n988), .A3(KEYINPUT118), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT118), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1070), .B(new_n1071), .C1(new_n1079), .C2(new_n1069), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n769), .A2(new_n251), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n773), .B1(new_n466), .B2(new_n215), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n756), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n841), .A2(G50), .B1(new_n809), .B2(new_n257), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n796), .A2(G77), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n382), .B1(new_n790), .B2(G143), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n792), .A2(new_n1005), .B1(new_n783), .B2(new_n812), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n202), .B2(new_n804), .C1(new_n399), .C2(new_n800), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n792), .A2(new_n1043), .B1(new_n783), .B2(new_n786), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n429), .B2(new_n800), .C1(new_n837), .C2(new_n804), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1040), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G294), .A2(new_n809), .B1(new_n790), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n287), .B1(new_n841), .B2(G303), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n468), .C2(new_n795), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1087), .A2(new_n1090), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1083), .B1(new_n1098), .B2(new_n772), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT119), .Z(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n762), .B2(new_n943), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1079), .B2(new_n755), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1080), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(G390));
  AOI21_X1  g0904(.A(new_n928), .B1(new_n880), .B2(new_n904), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n748), .A2(new_n695), .A3(new_n882), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1106), .A2(new_n883), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n891), .A2(new_n892), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n928), .B1(new_n921), .B2(new_n909), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n933), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n909), .A2(new_n738), .A3(new_n826), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1109), .B(new_n1112), .C1(new_n933), .C2(new_n1110), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n917), .A2(new_n658), .A3(new_n914), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n738), .A2(new_n826), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n921), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1112), .A2(new_n1118), .A3(new_n1107), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1114), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1071), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT120), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1122), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(KEYINPUT120), .A3(new_n1071), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1114), .A2(new_n755), .A3(new_n1115), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n757), .B1(new_n376), .B2(new_n831), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n382), .B1(new_n804), .B2(new_n399), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT121), .Z(new_n1135));
  AOI22_X1  g0935(.A1(G116), .A2(new_n816), .B1(new_n790), .B2(G294), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n466), .B2(new_n785), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1085), .B1(new_n429), .B2(new_n779), .C1(new_n837), .C2(new_n792), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n848), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n804), .A2(new_n1005), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n800), .A2(new_n207), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n287), .B1(new_n795), .B2(new_n812), .C1(new_n792), .C2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n783), .A2(new_n846), .B1(new_n785), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n779), .A2(new_n843), .B1(new_n789), .B2(new_n1147), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1135), .A2(new_n1139), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1133), .B1(new_n833), .B2(new_n1150), .C1(new_n933), .C2(new_n761), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1132), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1131), .A2(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n1116), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1123), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT123), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n912), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n934), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n894), .A2(KEYINPUT123), .A3(new_n910), .A4(G330), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n647), .B1(new_n314), .B2(new_n317), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n282), .A2(new_n692), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT122), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1163), .B(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n927), .B1(new_n930), .B2(new_n932), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n912), .B(new_n1157), .C1(new_n1168), .C2(new_n925), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1159), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1167), .B1(new_n1159), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1156), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1156), .B(KEYINPUT57), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1071), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n755), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n760), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n772), .A2(G50), .A3(new_n760), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n382), .B2(new_n302), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n612), .A2(new_n785), .B1(new_n837), .B2(new_n789), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n466), .A2(new_n779), .B1(new_n783), .B2(new_n429), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n302), .B(new_n382), .C1(new_n792), .C2(new_n468), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(new_n1001), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n801), .A2(G58), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1050), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n783), .A2(new_n1143), .B1(new_n785), .B2(new_n843), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n792), .A2(new_n1147), .B1(new_n779), .B2(new_n846), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G150), .C2(new_n796), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n804), .B2(new_n1145), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n801), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1190), .B1(new_n1189), .B2(new_n1188), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n757), .B(new_n1179), .C1(new_n1200), .C2(new_n772), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1178), .A2(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1177), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1176), .A2(new_n1203), .ZN(G375));
  NAND3_X1  g1004(.A1(new_n1120), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1128), .A2(new_n994), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n754), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1108), .A2(new_n760), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n290), .A2(new_n800), .B1(new_n804), .B2(new_n466), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n382), .B1(new_n789), .B2(new_n805), .C1(new_n612), .C2(new_n795), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n468), .A2(new_n779), .B1(new_n783), .B2(new_n837), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n792), .A2(new_n838), .B1(new_n785), .B2(new_n429), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT124), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n779), .A2(new_n1145), .B1(new_n785), .B2(new_n1005), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n287), .B1(new_n795), .B2(new_n207), .C1(new_n843), .C2(new_n783), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G132), .C2(new_n793), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n804), .A2(new_n812), .B1(new_n1143), .B2(new_n789), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT125), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT125), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1187), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n833), .B1(new_n1214), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n757), .B(new_n1222), .C1(new_n202), .C2(new_n831), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1207), .B1(new_n1208), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1206), .A2(new_n1224), .ZN(G381));
  NAND2_X1  g1025(.A1(new_n1177), .A2(new_n1202), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1062), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n1175), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1124), .A2(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1152), .B1(new_n1229), .B2(new_n1130), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n997), .A2(new_n1103), .A3(new_n1027), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n822), .B(new_n1061), .C1(new_n1064), .C2(new_n1067), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(G381), .A2(new_n1233), .A3(G384), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1228), .A2(new_n1230), .A3(new_n1232), .A4(new_n1234), .ZN(G407));
  NAND2_X1  g1035(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1236), .ZN(G409));
  NAND2_X1  g1037(.A1(new_n693), .A2(G213), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1156), .B(new_n994), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1230), .A2(new_n1203), .A3(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1205), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1120), .A2(new_n1116), .A3(KEYINPUT60), .A4(new_n1121), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1128), .A2(new_n1243), .A3(new_n1071), .A4(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1245), .B2(new_n1224), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(G384), .A3(new_n1224), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT62), .B1(new_n1241), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n693), .A2(G213), .A3(G2897), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1249), .B(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT61), .B1(new_n1241), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G375), .A2(G378), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1239), .A2(new_n1177), .A3(new_n1202), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1238), .B1(G378), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1249), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1254), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1250), .A2(new_n1253), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1103), .B1(new_n997), .B2(new_n1027), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1264), .A2(new_n1233), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1232), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1233), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(G390), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(new_n1231), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1262), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1265), .B1(new_n1232), .B2(new_n1263), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n1231), .A3(new_n1267), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1261), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1230), .B1(new_n1176), .B2(new_n1203), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1276), .A2(new_n1256), .A3(new_n1249), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT63), .B1(new_n1277), .B2(KEYINPUT126), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(new_n1241), .C2(new_n1249), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1253), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1275), .A2(new_n1283), .ZN(G405));
  AND3_X1   g1084(.A1(new_n1271), .A2(new_n1272), .A3(KEYINPUT127), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1259), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1254), .A2(new_n1236), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1270), .A2(new_n1273), .A3(new_n1249), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


