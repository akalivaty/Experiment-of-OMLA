//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT68), .B(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n472), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n479), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G138), .B1(new_n471), .B2(new_n472), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n487), .B2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n462), .A2(new_n470), .A3(new_n489), .A4(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n459), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n495), .A2(new_n499), .B1(new_n462), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n507), .A2(new_n508), .B1(G50), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n517), .B2(new_n511), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n504), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT72), .B1(new_n505), .B2(new_n506), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n514), .A2(new_n523), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n522), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(G51), .B2(new_n513), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n517), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n513), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n518), .A2(new_n521), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n518), .A2(G81), .A3(new_n521), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n513), .A2(G43), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n548), .A2(KEYINPUT73), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT73), .B1(new_n548), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  AOI22_X1  g133(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n506), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT74), .B1(new_n540), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n518), .A2(new_n563), .A3(G91), .A4(new_n521), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n513), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G74), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n506), .B1(new_n517), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(G49), .B2(new_n513), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n540), .B2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n504), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n506), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(KEYINPUT75), .B1(G48), .B2(new_n513), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n574), .A2(new_n575), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n506), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n518), .A2(G86), .A3(new_n521), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n513), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n540), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT76), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n506), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G54), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n519), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(new_n592), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n506), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n540), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n598), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n565), .A2(new_n567), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  XOR2_X1   g184(.A(KEYINPUT78), .B(G559), .Z(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(G860), .B2(new_n610), .ZN(G148));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n552), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n603), .A2(new_n610), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n462), .A2(new_n460), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(new_n624));
  AOI22_X1  g199(.A1(G123), .A2(new_n484), .B1(new_n480), .B2(G135), .ZN(new_n625));
  OAI221_X1 g200(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  OAI211_X1 g203(.A(new_n624), .B(new_n628), .C1(new_n622), .C2(new_n621), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(G14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(G401));
  XNOR2_X1  g220(.A(G2072), .B(G2078), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2084), .B(G2090), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT82), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n648), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n652), .B(new_n649), .C1(new_n646), .C2(new_n648), .ZN(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n654), .A2(new_n646), .A3(new_n648), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2096), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n664), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n668), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n665), .A2(KEYINPUT20), .A3(new_n668), .ZN(new_n673));
  OAI221_X1 g248(.A(new_n669), .B1(new_n668), .B2(new_n666), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT85), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n675), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NOR2_X1   g258(.A1(G168), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n683), .B2(G21), .ZN(new_n685));
  INV_X1    g260(.A(G1966), .ZN(new_n686));
  INV_X1    g261(.A(G2078), .ZN(new_n687));
  NAND2_X1  g262(.A1(G164), .A2(G29), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G27), .B2(G29), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT91), .B(KEYINPUT31), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G11), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT92), .B(G28), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n692), .B1(new_n694), .B2(new_n697), .C1(new_n627), .C2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G2084), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT24), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(G34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n477), .B2(G29), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n698), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n690), .B(new_n705), .C1(new_n699), .C2(new_n704), .ZN(new_n706));
  NOR2_X1   g281(.A1(G29), .A2(G35), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G162), .B2(G29), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2090), .ZN(new_n711));
  NOR2_X1   g286(.A1(G4), .A2(G16), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n603), .B2(G16), .ZN(new_n713));
  OAI22_X1  g288(.A1(new_n710), .A2(new_n711), .B1(G1348), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n689), .A2(new_n687), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n696), .A2(G33), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT25), .Z(new_n718));
  AOI22_X1  g293(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(new_n470), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n480), .A2(G139), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n696), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n715), .B1(new_n724), .B2(G2072), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n725), .B1(G2072), .B2(new_n724), .C1(new_n686), .C2(new_n685), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n706), .A2(new_n714), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n713), .A2(G1348), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n710), .A2(new_n711), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n696), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n484), .A2(G128), .ZN(new_n732));
  OAI221_X1 g307(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n480), .A2(G140), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n732), .A2(new_n733), .A3(new_n734), .A4(KEYINPUT89), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n731), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n683), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n683), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1961), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n460), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n484), .A2(G129), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT90), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G32), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n748), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n749), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n553), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G16), .B2(G19), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1341), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G1341), .B2(new_n762), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n683), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1956), .Z(new_n770));
  NOR3_X1   g345(.A1(new_n745), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G290), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT86), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n775));
  NAND2_X1  g350(.A1(G290), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n683), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G24), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n777), .A2(G1986), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(G1986), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(KEYINPUT87), .ZN(new_n782));
  AOI22_X1  g357(.A1(G119), .A2(new_n484), .B1(new_n480), .B2(G131), .ZN(new_n783));
  OAI221_X1 g358(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G25), .B(new_n785), .S(G29), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT35), .B(G1991), .Z(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n786), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(G166), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G16), .B2(G22), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  OR2_X1    g367(.A1(G6), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G305), .B2(new_n683), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  AOI22_X1  g370(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n792), .B2(new_n791), .ZN(new_n797));
  MUX2_X1   g372(.A(G23), .B(G288), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n794), .B2(new_n795), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n789), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n782), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n779), .A2(new_n807), .A3(new_n780), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT88), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n802), .B2(new_n803), .ZN(new_n810));
  OAI211_X1 g385(.A(KEYINPUT88), .B(KEYINPUT34), .C1(new_n797), .C2(new_n801), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n805), .A2(new_n806), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n812), .A2(new_n782), .A3(new_n804), .A4(new_n808), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT36), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n772), .B1(new_n813), .B2(new_n815), .ZN(G311));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n771), .ZN(G150));
  NAND2_X1  g393(.A1(new_n603), .A2(G559), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT38), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n513), .A2(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(new_n506), .B2(new_n822), .C1(new_n540), .C2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n552), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n552), .A2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n820), .B(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n829), .A2(new_n830), .A3(G860), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n824), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n833));
  XOR2_X1   g408(.A(new_n832), .B(new_n833), .Z(new_n834));
  OR2_X1    g409(.A1(new_n831), .A2(new_n834), .ZN(G145));
  AOI21_X1  g410(.A(new_n502), .B1(new_n737), .B2(new_n739), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n737), .A2(new_n502), .A3(new_n739), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n837), .A2(new_n754), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n754), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n722), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT96), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(new_n722), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n837), .A2(KEYINPUT95), .A3(new_n838), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT95), .B1(new_n837), .B2(new_n838), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n755), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n723), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n845), .A2(new_n846), .A3(new_n755), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n842), .B(new_n844), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n484), .A2(G130), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT97), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n470), .A2(G118), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(KEYINPUT98), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(KEYINPUT98), .B2(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n480), .A2(G142), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n852), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n785), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n620), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n627), .B(new_n477), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT100), .Z(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n850), .B2(new_n860), .ZN(new_n866));
  AOI21_X1  g441(.A(G37), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n850), .A2(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT99), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n850), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n861), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(KEYINPUT40), .B(new_n867), .C1(new_n872), .C2(new_n864), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n850), .A2(new_n870), .A3(new_n860), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n870), .B1(new_n850), .B2(new_n860), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n862), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n864), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT40), .B1(new_n879), .B2(new_n867), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n874), .A2(new_n880), .ZN(G395));
  NAND2_X1  g456(.A1(new_n827), .A2(new_n615), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n825), .A2(new_n614), .A3(new_n826), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n603), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n607), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n603), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT101), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n882), .A2(new_n888), .A3(new_n891), .A4(new_n883), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n886), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n897), .A2(new_n884), .A3(KEYINPUT102), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT102), .B1(new_n897), .B2(new_n884), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G288), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G305), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n893), .B(new_n907), .C1(new_n899), .C2(new_n898), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n902), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n902), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n824), .A2(new_n612), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(G295));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n912), .ZN(G331));
  NAND2_X1  g489(.A1(G301), .A2(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  NAND3_X1  g492(.A1(G301), .A2(KEYINPUT104), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(G168), .B1(KEYINPUT104), .B2(G301), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  AOI21_X1  g497(.A(G286), .B1(new_n922), .B2(G171), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n916), .A3(new_n918), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n921), .A2(new_n924), .A3(new_n826), .A4(new_n825), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(new_n889), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n924), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n827), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n928), .A3(new_n827), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n827), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n934), .A2(new_n925), .B1(new_n895), .B2(new_n896), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n936), .A3(new_n905), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n932), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n930), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n941), .B2(new_n927), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n905), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n942), .B2(new_n905), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n927), .A2(new_n934), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n940), .A2(new_n930), .A3(new_n926), .ZN(new_n947));
  INV_X1    g522(.A(new_n897), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n906), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n944), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n945), .A2(new_n950), .A3(KEYINPUT43), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n942), .A2(new_n905), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT43), .B1(new_n957), .B2(new_n945), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(G397));
  XNOR2_X1  g535(.A(new_n741), .B(G2067), .ZN(new_n961));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  INV_X1    g537(.A(new_n754), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT107), .B(G1384), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n502), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n468), .A2(new_n968), .A3(new_n475), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n970), .A2(KEYINPUT108), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(KEYINPUT108), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n964), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n785), .B(new_n787), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(G1996), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n755), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n980));
  OAI221_X1 g555(.A(new_n975), .B1(new_n973), .B2(new_n976), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1986), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n773), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT109), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n982), .B2(new_n773), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g562(.A1(G303), .A2(G8), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n491), .B2(new_n501), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n969), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g571(.A(KEYINPUT50), .B(G1384), .C1(new_n491), .C2(new_n501), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n969), .C1(KEYINPUT45), .C2(new_n994), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n998), .A2(new_n711), .B1(new_n1000), .B2(new_n792), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n992), .B(KEYINPUT111), .C1(new_n993), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n792), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n502), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n994), .A2(new_n995), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n711), .A3(new_n969), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n993), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n990), .A2(new_n991), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n994), .A2(new_n969), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n571), .B(G1976), .C1(new_n572), .C2(new_n540), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1014), .A2(G8), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(G8), .A3(new_n1016), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1015), .A2(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G305), .A2(G1981), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n577), .A2(new_n580), .A3(new_n1023), .A4(new_n581), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1002), .A2(new_n1012), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n969), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(new_n969), .C1(new_n994), .C2(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n686), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n998), .A2(new_n699), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(G8), .A3(G168), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n987), .B1(new_n1031), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT113), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT63), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n1044), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n987), .C1(new_n1031), .C2(new_n1041), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1050));
  OR2_X1    g625(.A1(G288), .A2(G1976), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1024), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1021), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1030), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1052), .A2(new_n1053), .B1(new_n1054), .B2(new_n1029), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n567), .B1(new_n565), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g633(.A(KEYINPUT117), .B(new_n560), .C1(new_n562), .C2(new_n564), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n607), .A2(KEYINPUT57), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT56), .B(G2072), .Z(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1000), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1032), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1064), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(KEYINPUT118), .A3(new_n999), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT114), .B(G1956), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n996), .B2(new_n997), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT115), .B(new_n1070), .C1(new_n996), .C2(new_n997), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1062), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n998), .A2(G1348), .B1(G2067), .B2(new_n1015), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n603), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1069), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n562), .A2(new_n564), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n1081), .B2(new_n560), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n565), .A2(new_n1057), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n567), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1084), .A2(new_n1056), .B1(KEYINPUT57), .B2(new_n607), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1077), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1073), .A2(new_n1074), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT121), .B1(new_n1088), .B2(new_n1062), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1089), .A2(KEYINPUT61), .B1(new_n1086), .B2(new_n1076), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n885), .C1(new_n1078), .C2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n603), .B(new_n1091), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1015), .A2(G2067), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1007), .A2(new_n969), .A3(new_n1008), .ZN(new_n1096));
  INV_X1    g671(.A(G1348), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1098), .A3(KEYINPUT60), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1078), .A2(new_n1092), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1093), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT45), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1006), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(new_n962), .A3(new_n969), .A4(new_n999), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1015), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1102), .B1(new_n1108), .B2(new_n553), .ZN(new_n1109));
  AOI211_X1 g684(.A(KEYINPUT120), .B(new_n552), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1110));
  NAND2_X1  g685(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1103), .B(new_n965), .C1(new_n491), .C2(new_n501), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1032), .A2(G1996), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1107), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n553), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT120), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1108), .A2(new_n1102), .A3(new_n553), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1111), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1101), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1090), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1089), .A2(KEYINPUT61), .A3(new_n1076), .A4(new_n1086), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1087), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1038), .A2(G168), .A3(new_n1039), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1037), .A2(new_n686), .B1(new_n699), .B2(new_n998), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(G168), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT51), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n993), .B1(new_n1127), .B2(G168), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1000), .B2(G2078), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT123), .B(G1961), .Z(new_n1136));
  NAND2_X1  g711(.A1(new_n1096), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n969), .A2(KEYINPUT53), .A3(new_n687), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n1138), .A2(new_n967), .A3(new_n1114), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(G171), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n687), .A2(KEYINPUT53), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1135), .B(new_n1137), .C1(new_n1037), .C2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1031), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1140), .A2(G171), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1144), .A2(G171), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT54), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g727(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1133), .B(new_n1147), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1049), .B(new_n1055), .C1(new_n1124), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1040), .A2(G286), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1131), .B1(new_n1130), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1126), .A2(KEYINPUT51), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT62), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1129), .A2(new_n1160), .A3(new_n1132), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1031), .A2(new_n1149), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT125), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1159), .A2(new_n1161), .A3(new_n1165), .A4(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n986), .B1(new_n1155), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n984), .A2(new_n973), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT46), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n977), .B(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n961), .A2(new_n963), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n973), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(KEYINPUT47), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(KEYINPUT47), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1170), .A2(new_n981), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n785), .A2(new_n788), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT126), .Z(new_n1179));
  OAI211_X1 g754(.A(new_n975), .B(new_n1179), .C1(new_n979), .C2(new_n980), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n742), .A2(G2067), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n973), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1168), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n879), .A2(new_n867), .ZN(new_n1186));
  INV_X1    g760(.A(G319), .ZN(new_n1187));
  OR2_X1    g761(.A1(G227), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g762(.A1(G401), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  OAI21_X1  g764(.A(new_n681), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1191), .B1(new_n1190), .B2(new_n1189), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n1186), .A2(new_n953), .A3(new_n1192), .ZN(G308));
  NAND3_X1  g767(.A1(new_n1186), .A2(new_n953), .A3(new_n1192), .ZN(G225));
endmodule


