//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(G58), .A2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n211), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n212), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G68), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n213), .A2(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(new_n202), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n214), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(KEYINPUT11), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT12), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n263), .B2(G68), .ZN(new_n264));
  INV_X1    g0064(.A(new_n263), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n250), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n205), .B2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n264), .B(new_n266), .C1(new_n268), .C2(new_n250), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n258), .B2(KEYINPUT11), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G226), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G97), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n273), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT65), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(new_n290), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n205), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n297), .A2(new_n283), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n295), .B1(G238), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n285), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(G169), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(G179), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n304), .B2(G169), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n271), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n301), .A2(G190), .A3(new_n303), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(G200), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n259), .A3(new_n270), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT72), .ZN(new_n315));
  INV_X1    g0115(.A(new_n249), .ZN(new_n316));
  INV_X1    g0116(.A(G159), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT66), .A2(G58), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT66), .A2(G58), .ZN(new_n320));
  OAI21_X1  g0120(.A(G68), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n217), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n322), .B2(G20), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n213), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n274), .A2(new_n206), .A3(new_n275), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT7), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n330), .A3(G68), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n323), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(new_n255), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n327), .B1(new_n326), .B2(new_n213), .ZN(new_n335));
  NOR4_X1   g0135(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT7), .A4(G20), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n335), .A2(new_n336), .A3(new_n250), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT66), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(KEYINPUT66), .A2(G58), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n216), .B1(new_n342), .B2(G68), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n343), .A2(new_n206), .B1(new_n317), .B2(new_n316), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n334), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(KEYINPUT8), .A3(new_n341), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT67), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n340), .A2(KEYINPUT67), .A3(KEYINPUT8), .A4(new_n341), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n339), .A2(KEYINPUT8), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AND4_X1   g0151(.A1(new_n263), .A2(new_n348), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n346), .B2(new_n347), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n267), .B1(new_n353), .B2(new_n349), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT73), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n268), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n263), .A3(new_n349), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n333), .A2(new_n345), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n235), .A2(G1698), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(G223), .B2(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT74), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n284), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n297), .A2(G232), .A3(new_n283), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n294), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(G179), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n283), .B1(new_n363), .B2(new_n366), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n294), .A2(new_n369), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT18), .B1(new_n361), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n345), .A2(new_n255), .A3(new_n332), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n355), .A2(new_n360), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n368), .A2(new_n370), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n372), .B2(new_n373), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n361), .B2(new_n387), .ZN(new_n388));
  AND4_X1   g0188(.A1(new_n382), .A2(new_n377), .A3(new_n378), .A4(new_n387), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n376), .B(new_n381), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT75), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(KEYINPUT75), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n252), .B1(new_n353), .B2(new_n349), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n249), .A2(G150), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n201), .B2(new_n206), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n255), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n263), .A2(G50), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(G50), .B2(new_n267), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT9), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n278), .A2(G222), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G223), .A2(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n276), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n284), .C1(G77), .C2(new_n276), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n298), .A2(G226), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n294), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n383), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(G200), .B2(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT10), .ZN(new_n411));
  INV_X1    g0211(.A(G169), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n400), .B(new_n413), .C1(G179), .C2(new_n407), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(new_n276), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n284), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n295), .B1(G244), .B2(new_n298), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n383), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(G200), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT15), .B(G87), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n252), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT8), .B(G58), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n202), .A2(new_n213), .B1(new_n426), .B2(new_n316), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n255), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n205), .A2(G20), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(new_n254), .A3(G77), .A4(new_n214), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n430), .B(KEYINPUT68), .Z(new_n431));
  NAND2_X1  g0231(.A1(new_n265), .A2(new_n202), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT69), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT69), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n428), .A2(new_n431), .A3(new_n435), .A4(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n423), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n422), .B1(new_n437), .B2(KEYINPUT70), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(KEYINPUT70), .B2(new_n437), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n421), .A2(new_n412), .ZN(new_n441));
  INV_X1    g0241(.A(G179), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n419), .A2(new_n420), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n411), .A2(new_n414), .A3(new_n439), .A4(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n315), .A2(new_n393), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n223), .A2(new_n280), .A3(new_n417), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT19), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n448), .A2(new_n273), .A3(new_n280), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT64), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G20), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n447), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n450), .A2(new_n452), .A3(G33), .A4(G97), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n448), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n276), .A2(new_n213), .A3(G68), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n255), .B1(new_n265), .B2(new_n424), .ZN(new_n459));
  INV_X1    g0259(.A(new_n255), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n205), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n263), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G87), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n224), .B1(new_n290), .B2(G1), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n205), .A2(new_n292), .A3(G45), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n283), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G238), .A2(G1698), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n222), .B2(G1698), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n470), .A2(new_n276), .B1(G33), .B2(G116), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n283), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G200), .ZN(new_n473));
  OAI211_X1 g0273(.A(G190), .B(new_n468), .C1(new_n471), .C2(new_n283), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n222), .A2(G1698), .ZN(new_n476));
  OAI221_X1 g0276(.A(new_n476), .B1(G238), .B2(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n283), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n468), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n412), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n442), .B(new_n468), .C1(new_n471), .C2(new_n283), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n424), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n463), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n459), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n465), .A2(new_n475), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n278), .A2(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n276), .A2(G244), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n326), .A2(new_n222), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n488), .B(new_n490), .C1(new_n491), .C2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n276), .A2(G250), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n278), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n284), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT5), .B1(new_n287), .B2(new_n289), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT5), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n205), .B(G45), .C1(new_n497), .C2(G41), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n283), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NOR4_X1   g0300(.A1(new_n496), .A2(new_n284), .A3(new_n498), .A4(new_n292), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n412), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT76), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n500), .B2(new_n501), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n287), .A2(new_n289), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n497), .ZN(new_n508));
  INV_X1    g0308(.A(new_n498), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(G274), .A3(new_n283), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n499), .A3(KEYINPUT76), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n506), .A2(new_n495), .A3(new_n442), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT6), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n513), .A2(new_n280), .A3(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(G97), .B(G107), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n516), .A2(new_n213), .B1(new_n202), .B2(new_n316), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n335), .A2(new_n336), .A3(new_n417), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n255), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n265), .A2(new_n280), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n463), .A2(G97), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n504), .A2(new_n512), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n506), .A2(new_n495), .A3(new_n511), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n520), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n515), .A2(new_n513), .ZN(new_n528));
  INV_X1    g0328(.A(new_n514), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n453), .B1(G77), .B2(new_n249), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT7), .B1(new_n453), .B2(new_n276), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(G107), .C1(KEYINPUT7), .C2(new_n329), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n527), .B1(new_n534), .B2(new_n255), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n383), .B2(new_n503), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n487), .B(new_n523), .C1(new_n526), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n525), .B(new_n535), .C1(new_n383), .C2(new_n503), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n523), .A4(new_n487), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n508), .A2(new_n509), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(G270), .A3(new_n283), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n278), .A2(G257), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G264), .A2(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n276), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n547), .B(new_n284), .C1(G303), .C2(new_n276), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n548), .A3(new_n510), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G169), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n254), .A2(new_n214), .B1(G20), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n488), .B1(new_n280), .B2(G33), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n453), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT20), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n263), .A2(G116), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n463), .B2(G116), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(KEYINPUT78), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT78), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n551), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n557), .A2(new_n559), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n557), .A2(KEYINPUT78), .A3(new_n559), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(KEYINPUT21), .A3(new_n551), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n544), .A2(new_n548), .A3(new_n510), .ZN(new_n571));
  OAI211_X1 g0371(.A(G179), .B(new_n571), .C1(new_n560), .C2(new_n561), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(G190), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n549), .A2(G200), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n567), .A2(new_n573), .A3(new_n568), .A4(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n564), .A2(new_n570), .A3(new_n572), .A4(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n276), .A2(new_n213), .A3(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n276), .A2(new_n213), .A3(new_n579), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT24), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n584), .C1(G20), .C2(new_n478), .ZN(new_n585));
  NOR2_X1   g0385(.A1(KEYINPUT23), .A2(G107), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n453), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n583), .A2(KEYINPUT24), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n460), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n581), .B(new_n587), .C1(new_n583), .C2(KEYINPUT24), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n262), .A2(G20), .A3(new_n417), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n593), .B(KEYINPUT80), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(KEYINPUT25), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(KEYINPUT25), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(G107), .B2(new_n463), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n599));
  OAI211_X1 g0399(.A(G250), .B(new_n278), .C1(new_n324), .C2(new_n325), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G294), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n284), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n543), .A2(G264), .A3(new_n283), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n510), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(G190), .A3(new_n510), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n592), .A2(new_n598), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT81), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n605), .A2(new_n610), .A3(G169), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n605), .B2(G169), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n605), .A2(new_n442), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n597), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n615), .A2(new_n595), .B1(new_n417), .B2(new_n462), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n591), .B2(new_n590), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n609), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n576), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n446), .A2(new_n542), .A3(new_n619), .ZN(G372));
  AOI21_X1  g0420(.A(new_n550), .B1(new_n567), .B2(new_n568), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n572), .B1(new_n621), .B2(KEYINPUT21), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n562), .A2(new_n563), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT82), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n614), .A2(new_n617), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT82), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n564), .A2(new_n570), .A3(new_n626), .A4(new_n572), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n609), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n537), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n459), .A2(new_n485), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n481), .A2(new_n482), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n487), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  OR3_X1    g0436(.A1(new_n635), .A2(new_n636), .A3(new_n523), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n635), .B2(new_n523), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n446), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n376), .A2(new_n381), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n444), .A2(KEYINPUT83), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n444), .A2(KEYINPUT83), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n313), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n310), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n388), .A2(new_n389), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n642), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n411), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n414), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n641), .A2(new_n652), .ZN(G369));
  NAND2_X1  g0453(.A1(new_n213), .A2(new_n262), .ZN(new_n654));
  OAI21_X1  g0454(.A(G213), .B1(new_n654), .B2(KEYINPUT27), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT84), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n655), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G343), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n567), .B2(new_n568), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n624), .B2(new_n627), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n576), .A2(new_n663), .ZN(new_n666));
  OR3_X1    g0466(.A1(new_n665), .A2(KEYINPUT85), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT86), .B(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT85), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT87), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT87), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n667), .A2(new_n673), .A3(new_n669), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n618), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n617), .B2(new_n662), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n625), .A2(new_n662), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n662), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n625), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n622), .A2(new_n623), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n681), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n209), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n507), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n205), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n447), .A2(G116), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n689), .A2(new_n690), .B1(new_n219), .B2(new_n688), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT28), .Z(new_n692));
  AOI21_X1  g0492(.A(new_n681), .B1(new_n631), .B2(new_n639), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n539), .A2(new_n523), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT88), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n683), .A2(new_n625), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n487), .A3(new_n609), .A4(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n681), .B1(new_n700), .B2(new_n639), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n695), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n542), .A2(new_n619), .A3(new_n662), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  INV_X1    g0504(.A(new_n472), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n607), .A2(new_n571), .A3(G179), .A4(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n706), .B2(new_n503), .ZN(new_n707));
  INV_X1    g0507(.A(new_n503), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n549), .A2(new_n442), .A3(new_n472), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT30), .A4(new_n607), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n571), .A2(G179), .A3(new_n705), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n524), .A3(new_n605), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n713), .B2(new_n681), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n703), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n702), .B1(new_n669), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n692), .B1(new_n718), .B2(G1), .ZN(G364));
  NAND2_X1  g0519(.A1(new_n667), .A2(new_n670), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n213), .A2(G13), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT89), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G45), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n689), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n214), .B1(G20), .B2(new_n412), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR4_X1   g0530(.A1(new_n213), .A2(new_n442), .A3(G190), .A4(new_n385), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n213), .A2(new_n442), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n732), .A2(new_n250), .B1(new_n202), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n385), .A2(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n453), .A2(new_n383), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n417), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n383), .A2(G179), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n213), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n280), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n737), .A2(G20), .A3(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G87), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n276), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n736), .A2(new_n739), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT32), .ZN(new_n748));
  NOR4_X1   g0548(.A1(new_n213), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(G159), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n733), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n385), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n750), .B1(G50), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n751), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n342), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n749), .A2(new_n748), .A3(G159), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n747), .A2(new_n753), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n749), .B(KEYINPUT91), .Z(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G329), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n276), .B1(new_n744), .B2(G303), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n761), .B2(new_n741), .ZN(new_n762));
  INV_X1    g0562(.A(new_n735), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(G311), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  INV_X1    g0565(.A(new_n738), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n731), .A2(new_n765), .B1(new_n766), .B2(G283), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G322), .A2(new_n754), .B1(new_n752), .B2(G326), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n759), .A2(new_n764), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n730), .B1(new_n757), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n244), .A2(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n687), .A2(new_n276), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(G45), .C2(new_n218), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n687), .A2(new_n326), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G355), .B1(new_n552), .B2(new_n687), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n723), .B(new_n729), .C1(new_n777), .C2(KEYINPUT90), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n777), .A2(KEYINPUT90), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n728), .B(new_n770), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n724), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT93), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n675), .ZN(new_n785));
  INV_X1    g0585(.A(new_n728), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n720), .B2(new_n668), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  INV_X1    g0590(.A(KEYINPUT94), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n439), .A2(new_n791), .A3(new_n444), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n681), .A2(new_n440), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n643), .B2(new_n644), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n439), .A2(KEYINPUT94), .A3(new_n444), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n792), .A2(new_n794), .B1(new_n795), .B2(new_n793), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n693), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n717), .A2(new_n669), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n786), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n758), .A2(G311), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n326), .B1(new_n743), .B2(new_n417), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n802), .B(new_n742), .C1(G283), .C2(new_n731), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n738), .A2(new_n223), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n763), .B2(G116), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G294), .A2(new_n754), .B1(new_n752), .B2(G303), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n801), .A2(new_n803), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n763), .A2(G159), .B1(G150), .B2(new_n731), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  INV_X1    g0609(.A(new_n752), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G143), .B2(new_n754), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n758), .A2(G132), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n766), .A2(G68), .ZN(new_n815));
  INV_X1    g0615(.A(new_n741), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n342), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n326), .B1(new_n744), .B2(G50), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n814), .A2(new_n815), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n807), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n729), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n729), .A2(new_n721), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n728), .B1(new_n202), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n821), .B(new_n823), .C1(new_n796), .C2(new_n722), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n800), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  OR2_X1    g0626(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n827), .A2(G116), .A3(new_n215), .A4(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n830));
  XNOR2_X1  g0630(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n219), .A2(G77), .A3(new_n321), .ZN(new_n832));
  INV_X1    g0632(.A(G50), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(KEYINPUT96), .B1(new_n833), .B2(G68), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(KEYINPUT96), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n205), .A2(G13), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT99), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n377), .A2(new_n378), .A3(new_n387), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n379), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n377), .A2(new_n378), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n661), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n843), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n838), .A2(new_n844), .B1(new_n390), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n375), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n377), .A2(new_n378), .A3(new_n387), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n850), .B2(new_n845), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n843), .A3(new_n839), .A4(new_n849), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(KEYINPUT99), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n323), .A2(new_n331), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n334), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n333), .A2(new_n856), .B1(new_n355), .B2(new_n360), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n660), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n390), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n857), .B2(new_n375), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n860), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n852), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT100), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n390), .A2(new_n845), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n844), .A2(new_n838), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n853), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT100), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n390), .A2(new_n858), .B1(new_n861), .B2(new_n852), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT39), .B1(new_n873), .B2(KEYINPUT38), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(new_n863), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n866), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n866), .A2(new_n875), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n310), .A2(new_n681), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n681), .A2(new_n444), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n693), .B2(new_n796), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n662), .B1(new_n259), .B2(new_n270), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n308), .B2(new_n309), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT97), .ZN(new_n891));
  INV_X1    g0691(.A(new_n889), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n310), .A2(new_n313), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT97), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n889), .B(new_n894), .C1(new_n308), .C2(new_n309), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n888), .A2(KEYINPUT98), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT98), .B1(new_n888), .B2(new_n897), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n898), .B(new_n899), .C1(new_n877), .C2(new_n876), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n642), .A2(new_n660), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n886), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n651), .B1(new_n702), .B2(new_n446), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n902), .B(new_n903), .Z(new_n904));
  NAND4_X1  g0704(.A1(new_n717), .A2(new_n796), .A3(KEYINPUT40), .A4(new_n896), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n871), .A2(new_n863), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(KEYINPUT102), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT102), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n854), .A2(new_n877), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(new_n905), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n717), .A2(new_n796), .A3(new_n896), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n876), .A2(new_n877), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n446), .A2(new_n717), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n668), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n904), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n205), .B2(new_n726), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n904), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n837), .B1(new_n923), .B2(new_n924), .ZN(G367));
  NOR2_X1   g0725(.A1(new_n723), .A2(new_n729), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n209), .B2(new_n424), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n772), .B2(new_n240), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n728), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n723), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n662), .A2(new_n465), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n634), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n635), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n738), .A2(new_n280), .ZN(new_n934));
  INV_X1    g0734(.A(G283), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n732), .A2(new_n761), .B1(new_n935), .B2(new_n735), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n934), .B(new_n936), .C1(G317), .C2(new_n749), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n743), .A2(new_n552), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT46), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n276), .B(new_n939), .C1(G107), .C2(new_n816), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n752), .A2(G311), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n754), .A2(G303), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n937), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n738), .A2(new_n202), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n749), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n945), .B1(new_n732), .B2(new_n317), .C1(new_n809), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n816), .A2(G68), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n326), .B1(new_n744), .B2(new_n342), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G50), .B2(new_n763), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n754), .A2(G150), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n752), .A2(G143), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n943), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  OAI221_X1 g0756(.A(new_n929), .B1(new_n930), .B2(new_n933), .C1(new_n956), .C2(new_n730), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n684), .A2(new_n676), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n681), .A2(new_n522), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n698), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n662), .A2(new_n523), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n523), .B1(new_n961), .B2(new_n625), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n662), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT103), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n964), .A2(new_n966), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n933), .B(KEYINPUT43), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n679), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n672), .B2(new_n674), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n961), .A2(new_n962), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n974), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n727), .A2(G1), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT105), .ZN(new_n982));
  INV_X1    g0782(.A(new_n718), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n959), .B1(new_n679), .B2(new_n684), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n675), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n984), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n672), .B2(new_n674), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n718), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n685), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT44), .B1(new_n977), .B2(new_n685), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n977), .A2(KEYINPUT45), .A3(new_n685), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT45), .B1(new_n977), .B2(new_n685), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n989), .B(new_n990), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n976), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n993), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(new_n680), .A3(KEYINPUT104), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT104), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n976), .B2(new_n993), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n983), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n688), .B(KEYINPUT41), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n982), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n958), .B1(new_n980), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n772), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n237), .A2(G45), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT106), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n426), .A2(G50), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n690), .ZN(new_n1012));
  AOI211_X1 g0812(.A(G45), .B(new_n1012), .C1(G68), .C2(G77), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1007), .B(new_n1009), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n774), .A2(new_n1012), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(G107), .B2(new_n209), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n926), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G50), .A2(new_n754), .B1(new_n752), .B2(G159), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n816), .A2(new_n484), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n744), .A2(G77), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n276), .A3(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n934), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n356), .A2(new_n731), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT107), .B(G150), .Z(new_n1024));
  AOI22_X1  g0824(.A1(new_n763), .A2(G68), .B1(new_n749), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1018), .A2(new_n1022), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n276), .B1(new_n749), .B2(G326), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n741), .A2(new_n935), .B1(new_n761), .B2(new_n743), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n763), .A2(G303), .B1(G311), .B2(new_n731), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n754), .A2(G317), .ZN(new_n1030));
  INV_X1    g0830(.A(G322), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1030), .C1(new_n1031), .C2(new_n810), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1027), .B1(new_n552), .B2(new_n738), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1026), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n729), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1017), .A2(new_n786), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n975), .B2(new_n723), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n985), .A2(new_n987), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n982), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1043), .A2(new_n718), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n988), .A2(new_n688), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  XOR2_X1   g0848(.A(new_n994), .B(KEYINPUT108), .Z(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n1001), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n988), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n688), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n996), .B2(new_n1001), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(new_n1001), .A3(new_n1044), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n926), .B1(new_n280), .B2(new_n209), .C1(new_n1007), .C2(new_n247), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n786), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n816), .A2(G77), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n735), .B2(new_n426), .C1(new_n732), .C2(new_n833), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT111), .Z(new_n1060));
  AOI22_X1  g0860(.A1(G150), .A2(new_n752), .B1(new_n754), .B2(G159), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n749), .A2(G143), .B1(G68), .B2(new_n744), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT110), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT110), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n326), .B(new_n804), .C1(new_n1064), .C2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1060), .A2(new_n1063), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G311), .A2(new_n754), .B1(new_n752), .B2(G317), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT112), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  AOI22_X1  g0872(.A1(new_n763), .A2(G294), .B1(G303), .B2(new_n731), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1031), .B2(new_n946), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n326), .B1(new_n935), .B2(new_n743), .C1(new_n741), .C2(new_n552), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1074), .A2(new_n739), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1069), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1057), .B1(new_n1077), .B2(new_n729), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n977), .B2(new_n930), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1054), .A2(new_n1055), .A3(new_n1079), .ZN(G390));
  NOR2_X1   g0880(.A1(new_n393), .A2(new_n445), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n315), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1081), .A2(new_n1082), .A3(G330), .A4(new_n717), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n446), .A2(new_n1085), .A3(G330), .A4(new_n717), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n887), .B1(new_n701), .B2(new_n796), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n717), .A2(G330), .A3(new_n796), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n896), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n796), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n798), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n896), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1095), .A3(new_n896), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1089), .A2(new_n896), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n897), .B1(new_n798), .B2(new_n1091), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n888), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n903), .B(new_n1087), .C1(new_n1097), .C2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n884), .B1(new_n888), .B2(new_n897), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n880), .A2(new_n882), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n884), .B(new_n907), .C1(new_n1088), .C2(new_n897), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT113), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(KEYINPUT113), .B(new_n1098), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1102), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1098), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1087), .A2(new_n903), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1090), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1105), .A2(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1100), .A2(new_n888), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .A4(new_n1107), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1112), .A2(new_n1123), .A3(new_n688), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1116), .A2(new_n1044), .A3(new_n1122), .A4(new_n1107), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n822), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n758), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n761), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n815), .A2(new_n1058), .A3(new_n326), .A4(new_n745), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n732), .A2(new_n417), .B1(new_n280), .B2(new_n735), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n754), .A2(G116), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n810), .B2(new_n935), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n276), .B1(new_n738), .B2(new_n833), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n758), .B2(G125), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT117), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n744), .A2(new_n1024), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT53), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G128), .A2(new_n752), .B1(new_n754), .B2(G132), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(KEYINPUT53), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G159), .B2(new_n816), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT54), .B(G143), .Z(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT116), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1143), .A2(new_n763), .B1(G137), .B2(new_n731), .ZN(new_n1144));
  AND4_X1   g0944(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1133), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n786), .B1(new_n356), .B2(new_n1126), .C1(new_n1146), .C2(new_n730), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT118), .Z(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n883), .B2(new_n722), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1125), .A2(KEYINPUT119), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT119), .B1(new_n1125), .B2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1124), .B1(new_n1150), .B2(new_n1151), .ZN(G378));
  AOI21_X1  g0952(.A(KEYINPUT102), .B1(new_n906), .B2(new_n907), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n910), .A2(new_n905), .A3(new_n909), .ZN(new_n1154));
  OAI211_X1 g0954(.A(G330), .B(new_n916), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n411), .A2(new_n414), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n661), .A2(new_n400), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n912), .A2(new_n1160), .A3(G330), .A4(new_n916), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n902), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n883), .A2(new_n885), .B1(new_n642), .B2(new_n660), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1166), .A2(new_n1162), .A3(new_n900), .A4(new_n1163), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1044), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n786), .B1(G50), .B2(new_n1126), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n276), .A2(new_n507), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G50), .B(new_n1171), .C1(new_n273), .C2(new_n286), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n738), .B1(new_n340), .B2(new_n341), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n731), .A2(G97), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(new_n948), .A3(new_n1020), .A4(new_n1171), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(new_n484), .C2(new_n763), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G107), .A2(new_n754), .B1(new_n752), .B2(G116), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n935), .C2(new_n1127), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1172), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n752), .A2(G125), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n816), .A2(G150), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1143), .A2(new_n744), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n763), .A2(G137), .B1(G132), .B2(new_n731), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G128), .C2(new_n754), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n766), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n749), .C2(G124), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1180), .B1(new_n1179), .B2(new_n1178), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1170), .B1(new_n1194), .B2(new_n729), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1160), .B2(new_n722), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1169), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1110), .A2(new_n1102), .A3(new_n1111), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n1201), .B2(new_n1117), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(KEYINPUT121), .B(new_n1200), .C1(new_n1201), .C2(new_n1117), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1117), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1123), .A2(new_n1207), .B1(new_n1167), .B2(new_n1165), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n688), .B1(new_n1208), .B2(KEYINPUT57), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1198), .B1(new_n1206), .B2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n897), .A2(new_n721), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n786), .B1(G68), .B2(new_n1126), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n758), .A2(G303), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n276), .B1(new_n744), .B2(G97), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n945), .A2(new_n1019), .A3(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n763), .A2(G107), .B1(G116), .B2(new_n731), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G283), .A2(new_n754), .B1(new_n752), .B2(G294), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n758), .A2(G128), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n276), .B1(new_n743), .B2(new_n317), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1221), .B(new_n1173), .C1(G50), .C2(new_n816), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n754), .A2(G137), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n731), .A2(new_n1143), .B1(new_n763), .B2(G150), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n752), .A2(G132), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT122), .Z(new_n1227));
  OAI21_X1  g1027(.A(new_n1219), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1213), .B1(new_n1228), .B2(new_n729), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1211), .A2(new_n1044), .B1(new_n1212), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1003), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1102), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1211), .A2(new_n1207), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  INV_X1    g1034(.A(new_n1205), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1123), .A2(new_n1207), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT121), .B1(new_n1236), .B2(new_n1200), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1168), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1052), .B1(new_n1239), .B2(new_n1199), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1197), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n1005), .A4(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G343), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G213), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1241), .A2(new_n1244), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  OAI211_X1 g1050(.A(G378), .B(new_n1198), .C1(new_n1206), .C2(new_n1209), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1197), .B1(new_n1208), .B2(new_n1231), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(G378), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1233), .A2(KEYINPUT60), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1233), .A2(KEYINPUT60), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1121), .A2(new_n1052), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G384), .A3(new_n1230), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1258), .B2(new_n1230), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1254), .A2(new_n1247), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1258), .A2(new_n1230), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n825), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1248), .A2(G2897), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1259), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(new_n1266), .B2(new_n1259), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1252), .A2(G378), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1241), .B2(G378), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1273), .B2(new_n1248), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1248), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1262), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1264), .A2(new_n1274), .A3(new_n1275), .A4(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(G396), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1005), .B2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(new_n789), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n980), .A2(new_n1004), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n958), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G390), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1282), .A2(new_n1285), .A3(G390), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1279), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(KEYINPUT123), .B(new_n1271), .C1(new_n1273), .C2(new_n1248), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT123), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G2897), .B(new_n1248), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1268), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1293), .B1(new_n1276), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1282), .A2(new_n1285), .A3(G390), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1275), .B1(new_n1298), .B2(new_n1286), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1263), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT125), .B1(new_n1263), .B2(new_n1300), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1276), .A2(new_n1303), .A3(KEYINPUT63), .A4(new_n1262), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1297), .A2(new_n1301), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1291), .A2(new_n1305), .ZN(G405));
  NOR2_X1   g1106(.A1(new_n1241), .A2(G378), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1251), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1262), .B(KEYINPUT126), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1289), .A2(KEYINPUT127), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1289), .A2(KEYINPUT127), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1262), .A2(KEYINPUT126), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1307), .A2(new_n1308), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .A4(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1318));
  OAI211_X1 g1118(.A(KEYINPUT127), .B(new_n1289), .C1(new_n1318), .C2(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(G402));
endmodule


