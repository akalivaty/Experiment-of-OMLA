

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783;

  XNOR2_X1 U373 ( .A(G143), .B(G122), .ZN(n591) );
  XNOR2_X1 U374 ( .A(G128), .B(G110), .ZN(n531) );
  XOR2_X2 U375 ( .A(n450), .B(n518), .Z(n412) );
  XOR2_X2 U376 ( .A(n530), .B(n529), .Z(n411) );
  XOR2_X2 U377 ( .A(KEYINPUT75), .B(KEYINPUT34), .Z(n618) );
  XNOR2_X1 U378 ( .A(G116), .B(G146), .ZN(n524) );
  BUF_X1 U379 ( .A(G113), .Z(n466) );
  XOR2_X1 U380 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n352) );
  AND2_X1 U381 ( .A1(n379), .A2(n493), .ZN(n353) );
  AND2_X2 U382 ( .A1(n361), .A2(n363), .ZN(n360) );
  NOR2_X1 U383 ( .A1(G902), .A2(n749), .ZN(n546) );
  NOR2_X1 U384 ( .A1(n741), .A2(G902), .ZN(n559) );
  INV_X1 U385 ( .A(n565), .ZN(n536) );
  INV_X4 U386 ( .A(G128), .ZN(n494) );
  NAND2_X1 U387 ( .A1(n370), .A2(n513), .ZN(n443) );
  OR2_X1 U388 ( .A1(n375), .A2(G902), .ZN(n391) );
  INV_X1 U389 ( .A(n354), .ZN(n398) );
  INV_X1 U390 ( .A(n572), .ZN(n354) );
  OR2_X1 U391 ( .A1(G237), .A2(G902), .ZN(n573) );
  INV_X1 U392 ( .A(KEYINPUT44), .ZN(n369) );
  INV_X1 U393 ( .A(KEYINPUT85), .ZN(n384) );
  INV_X1 U394 ( .A(KEYINPUT3), .ZN(n527) );
  INV_X1 U395 ( .A(KEYINPUT91), .ZN(n505) );
  INV_X1 U396 ( .A(KEYINPUT30), .ZN(n377) );
  XOR2_X1 U397 ( .A(G140), .B(G137), .Z(n548) );
  INV_X1 U398 ( .A(KEYINPUT6), .ZN(n390) );
  OR2_X1 U399 ( .A1(n675), .A2(n697), .ZN(n403) );
  NAND2_X1 U400 ( .A1(n372), .A2(n471), .ZN(n697) );
  INV_X1 U401 ( .A(n374), .ZN(n372) );
  AND2_X1 U402 ( .A1(n357), .A2(n389), .ZN(n356) );
  NOR2_X1 U403 ( .A1(n671), .A2(n693), .ZN(n421) );
  AND2_X1 U404 ( .A1(n444), .A2(n443), .ZN(n408) );
  NAND2_X1 U405 ( .A1(n380), .A2(n381), .ZN(n357) );
  XNOR2_X1 U406 ( .A(n389), .B(G101), .ZN(G3) );
  NAND2_X1 U407 ( .A1(n366), .A2(n487), .ZN(n359) );
  NAND2_X1 U408 ( .A1(n668), .A2(n480), .ZN(n669) );
  NAND2_X1 U409 ( .A1(n370), .A2(n451), .ZN(n389) );
  XNOR2_X1 U410 ( .A(n656), .B(KEYINPUT40), .ZN(n371) );
  XNOR2_X1 U411 ( .A(n628), .B(n352), .ZN(n382) );
  AND2_X1 U412 ( .A1(n430), .A2(n405), .ZN(n686) );
  AND2_X1 U413 ( .A1(n482), .A2(n404), .ZN(n405) );
  XNOR2_X1 U414 ( .A(n499), .B(n498), .ZN(n781) );
  NOR2_X1 U415 ( .A1(n653), .A2(n661), .ZN(n655) );
  INV_X1 U416 ( .A(n688), .ZN(n394) );
  INV_X1 U417 ( .A(n691), .ZN(n395) );
  NOR2_X1 U418 ( .A1(n650), .A2(n715), .ZN(n386) );
  INV_X1 U419 ( .A(n720), .ZN(n396) );
  AND2_X1 U420 ( .A1(n493), .A2(n384), .ZN(n362) );
  INV_X1 U421 ( .A(n662), .ZN(n501) );
  AND2_X1 U422 ( .A1(n502), .A2(n492), .ZN(n491) );
  AND2_X1 U423 ( .A1(n614), .A2(n646), .ZN(n610) );
  AND2_X1 U424 ( .A1(n644), .A2(n452), .ZN(n513) );
  XNOR2_X1 U425 ( .A(n378), .B(n377), .ZN(n376) );
  NAND2_X1 U426 ( .A1(n649), .A2(n700), .ZN(n378) );
  NOR2_X1 U427 ( .A1(n452), .A2(n637), .ZN(n451) );
  XNOR2_X1 U428 ( .A(n715), .B(n390), .ZN(n637) );
  NAND2_X1 U429 ( .A1(n710), .A2(n614), .ZN(n712) );
  XNOR2_X1 U430 ( .A(n715), .B(KEYINPUT106), .ZN(n649) );
  INV_X1 U431 ( .A(n439), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n483), .B(n767), .ZN(n741) );
  NAND2_X1 U433 ( .A1(n673), .A2(KEYINPUT65), .ZN(n439) );
  XNOR2_X1 U434 ( .A(n547), .B(n548), .ZN(n767) );
  XNOR2_X1 U435 ( .A(n608), .B(n406), .ZN(n547) );
  XNOR2_X1 U436 ( .A(n554), .B(n553), .ZN(n753) );
  XNOR2_X1 U437 ( .A(n566), .B(n528), .ZN(n608) );
  XNOR2_X1 U438 ( .A(n555), .B(KEYINPUT74), .ZN(n556) );
  XNOR2_X1 U439 ( .A(n505), .B(KEYINPUT72), .ZN(n504) );
  XOR2_X2 U440 ( .A(G122), .B(G116), .Z(n604) );
  XOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n569) );
  XNOR2_X2 U442 ( .A(G104), .B(G110), .ZN(n552) );
  XNOR2_X1 U443 ( .A(G107), .B(KEYINPUT90), .ZN(n553) );
  NAND2_X1 U444 ( .A1(n382), .A2(n385), .ZN(n380) );
  AND2_X1 U445 ( .A1(n613), .A2(n615), .ZN(n370) );
  XNOR2_X1 U446 ( .A(n355), .B(n467), .ZN(n449) );
  NAND2_X1 U447 ( .A1(n358), .A2(n356), .ZN(n355) );
  NAND2_X1 U448 ( .A1(n360), .A2(n359), .ZN(n358) );
  NAND2_X1 U449 ( .A1(n364), .A2(n453), .ZN(n361) );
  AND2_X1 U450 ( .A1(n379), .A2(n362), .ZN(n366) );
  NAND2_X1 U451 ( .A1(n365), .A2(n383), .ZN(n363) );
  NAND2_X1 U452 ( .A1(n379), .A2(n455), .ZN(n364) );
  NAND2_X1 U453 ( .A1(n365), .A2(n491), .ZN(n487) );
  INV_X1 U454 ( .A(n620), .ZN(n365) );
  NOR2_X1 U455 ( .A1(n367), .A2(n439), .ZN(n438) );
  NAND2_X1 U456 ( .A1(n433), .A2(n367), .ZN(n432) );
  XNOR2_X2 U457 ( .A(n630), .B(n629), .ZN(n367) );
  NAND2_X1 U458 ( .A1(n368), .A2(KEYINPUT44), .ZN(n446) );
  INV_X1 U459 ( .A(n443), .ZN(n368) );
  AND2_X1 U460 ( .A1(n443), .A2(n369), .ZN(n445) );
  XNOR2_X1 U461 ( .A(n443), .B(G110), .ZN(G12) );
  NAND2_X1 U462 ( .A1(n371), .A2(n783), .ZN(n418) );
  XNOR2_X1 U463 ( .A(n371), .B(G131), .ZN(G33) );
  NAND2_X1 U464 ( .A1(n497), .A2(n495), .ZN(n374) );
  NAND2_X1 U465 ( .A1(n374), .A2(n373), .ZN(n437) );
  NOR2_X1 U466 ( .A1(n374), .A2(KEYINPUT65), .ZN(n433) );
  XNOR2_X1 U467 ( .A(n374), .B(n769), .ZN(n771) );
  XNOR2_X1 U468 ( .A(n375), .B(KEYINPUT110), .ZN(n529) );
  XNOR2_X1 U469 ( .A(n423), .B(n422), .ZN(n375) );
  NAND2_X1 U470 ( .A1(n652), .A2(n376), .ZN(n661) );
  NAND2_X2 U471 ( .A1(n620), .A2(KEYINPUT35), .ZN(n379) );
  INV_X1 U472 ( .A(n667), .ZN(n381) );
  OR2_X1 U473 ( .A1(n382), .A2(n394), .ZN(n689) );
  OR2_X1 U474 ( .A1(n382), .A2(n395), .ZN(n692) );
  AND2_X1 U475 ( .A1(n491), .A2(n489), .ZN(n383) );
  XNOR2_X2 U476 ( .A(n619), .B(n618), .ZN(n620) );
  BUF_X2 U477 ( .A(n456), .Z(n402) );
  INV_X1 U478 ( .A(n385), .ZN(n678) );
  NAND2_X1 U479 ( .A1(n617), .A2(n386), .ZN(n385) );
  XNOR2_X2 U480 ( .A(n388), .B(n387), .ZN(n613) );
  INV_X1 U481 ( .A(n611), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n617), .A2(n610), .ZN(n388) );
  NAND2_X1 U483 ( .A1(n627), .A2(n637), .ZN(n616) );
  XNOR2_X2 U484 ( .A(n391), .B(G472), .ZN(n715) );
  XNOR2_X2 U485 ( .A(n392), .B(n574), .ZN(n658) );
  NAND2_X1 U486 ( .A1(n631), .A2(n700), .ZN(n392) );
  XNOR2_X2 U487 ( .A(n393), .B(n520), .ZN(n631) );
  NAND2_X1 U488 ( .A1(n397), .A2(n398), .ZN(n393) );
  AND2_X1 U489 ( .A1(n617), .A2(n396), .ZN(n628) );
  XNOR2_X2 U490 ( .A(n582), .B(KEYINPUT0), .ZN(n617) );
  XNOR2_X1 U491 ( .A(n464), .B(n399), .ZN(n397) );
  INV_X1 U492 ( .A(n400), .ZN(n399) );
  INV_X1 U493 ( .A(n516), .ZN(n400) );
  XNOR2_X2 U494 ( .A(n752), .B(n567), .ZN(n464) );
  BUF_X1 U495 ( .A(n564), .Z(n401) );
  INV_X1 U496 ( .A(n779), .ZN(n444) );
  INV_X1 U497 ( .A(G134), .ZN(n528) );
  OR2_X1 U498 ( .A1(n673), .A2(KEYINPUT65), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n686), .B(n481), .ZN(n480) );
  INV_X1 U500 ( .A(KEYINPUT47), .ZN(n481) );
  NAND2_X1 U501 ( .A1(n408), .A2(n778), .ZN(n440) );
  NAND2_X1 U502 ( .A1(n407), .A2(n442), .ZN(n441) );
  INV_X1 U503 ( .A(n651), .ZN(n477) );
  INV_X1 U504 ( .A(KEYINPUT15), .ZN(n478) );
  XNOR2_X1 U505 ( .A(KEYINPUT89), .B(G902), .ZN(n479) );
  XNOR2_X1 U506 ( .A(n526), .B(n522), .ZN(n424) );
  XNOR2_X1 U507 ( .A(n421), .B(n420), .ZN(n419) );
  XNOR2_X1 U508 ( .A(n418), .B(n409), .ZN(n417) );
  INV_X1 U509 ( .A(KEYINPUT69), .ZN(n420) );
  NAND2_X1 U510 ( .A1(n663), .A2(KEYINPUT35), .ZN(n493) );
  INV_X1 U511 ( .A(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U512 ( .A(n602), .B(n469), .ZN(n606) );
  NOR2_X1 U513 ( .A1(n438), .A2(n435), .ZN(n434) );
  NAND2_X1 U514 ( .A1(n427), .A2(n425), .ZN(n430) );
  XNOR2_X1 U515 ( .A(n567), .B(n465), .ZN(n483) );
  XNOR2_X1 U516 ( .A(n551), .B(n557), .ZN(n465) );
  NOR2_X1 U517 ( .A1(n621), .A2(n490), .ZN(n489) );
  XOR2_X1 U518 ( .A(KEYINPUT76), .B(G137), .Z(n525) );
  INV_X1 U519 ( .A(KEYINPUT84), .ZN(n467) );
  NOR2_X1 U520 ( .A1(G953), .A2(G237), .ZN(n588) );
  XNOR2_X1 U521 ( .A(n603), .B(n470), .ZN(n469) );
  INV_X1 U522 ( .A(KEYINPUT104), .ZN(n470) );
  XOR2_X1 U523 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n603) );
  XOR2_X1 U524 ( .A(G140), .B(G131), .Z(n594) );
  XNOR2_X1 U525 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n585) );
  XOR2_X1 U526 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n586) );
  INV_X1 U527 ( .A(KEYINPUT82), .ZN(n629) );
  INV_X1 U528 ( .A(KEYINPUT70), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n709), .A2(n477), .ZN(n476) );
  NOR2_X1 U530 ( .A1(n644), .A2(n431), .ZN(n426) );
  XNOR2_X1 U531 ( .A(n523), .B(n401), .ZN(n422) );
  XNOR2_X1 U532 ( .A(n547), .B(n424), .ZN(n423) );
  NOR2_X1 U533 ( .A1(n696), .A2(n496), .ZN(n495) );
  INV_X1 U534 ( .A(n695), .ZN(n496) );
  XNOR2_X1 U535 ( .A(n604), .B(KEYINPUT16), .ZN(n563) );
  XNOR2_X1 U536 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U537 ( .A(n566), .B(n565), .ZN(n517) );
  AND2_X1 U538 ( .A1(n430), .A2(n404), .ZN(n666) );
  NAND2_X1 U539 ( .A1(n487), .A2(n353), .ZN(n778) );
  INV_X1 U540 ( .A(KEYINPUT32), .ZN(n514) );
  INV_X1 U541 ( .A(n473), .ZN(n482) );
  INV_X1 U542 ( .A(KEYINPUT107), .ZN(n498) );
  NOR2_X1 U543 ( .A1(n661), .A2(n500), .ZN(n499) );
  NAND2_X1 U544 ( .A1(n502), .A2(n501), .ZN(n500) );
  INV_X1 U545 ( .A(KEYINPUT122), .ZN(n508) );
  INV_X1 U546 ( .A(KEYINPUT60), .ZN(n458) );
  XNOR2_X1 U547 ( .A(n739), .B(n468), .ZN(n742) );
  XNOR2_X1 U548 ( .A(n741), .B(n740), .ZN(n468) );
  XNOR2_X1 U549 ( .A(n479), .B(n478), .ZN(n572) );
  XNOR2_X1 U550 ( .A(KEYINPUT108), .B(n645), .ZN(n404) );
  INV_X1 U551 ( .A(n663), .ZN(n502) );
  XNOR2_X1 U552 ( .A(n571), .B(n517), .ZN(n516) );
  XOR2_X1 U553 ( .A(KEYINPUT4), .B(G131), .Z(n406) );
  AND2_X1 U554 ( .A1(n447), .A2(n446), .ZN(n407) );
  INV_X1 U555 ( .A(n649), .ZN(n644) );
  XOR2_X1 U556 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n409) );
  XOR2_X1 U557 ( .A(n744), .B(n743), .Z(n410) );
  XOR2_X1 U558 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n413) );
  XNOR2_X1 U559 ( .A(KEYINPUT88), .B(n521), .ZN(n751) );
  INV_X1 U560 ( .A(n751), .ZN(n462) );
  XNOR2_X1 U561 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n414) );
  XOR2_X1 U562 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n415) );
  XNOR2_X1 U563 ( .A(n416), .B(n413), .ZN(n497) );
  NAND2_X1 U564 ( .A1(n419), .A2(n417), .ZN(n416) );
  NAND2_X1 U565 ( .A1(n429), .A2(n426), .ZN(n425) );
  NAND2_X1 U566 ( .A1(n428), .A2(n431), .ZN(n427) );
  NAND2_X1 U567 ( .A1(n429), .A2(n649), .ZN(n428) );
  INV_X1 U568 ( .A(n643), .ZN(n429) );
  INV_X1 U569 ( .A(KEYINPUT28), .ZN(n431) );
  NAND2_X1 U570 ( .A1(n434), .A2(n432), .ZN(n457) );
  NAND2_X1 U571 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U572 ( .A1(n441), .A2(n440), .ZN(n448) );
  NAND2_X1 U573 ( .A1(n445), .A2(n444), .ZN(n442) );
  NAND2_X1 U574 ( .A1(n779), .A2(KEYINPUT44), .ZN(n447) );
  NAND2_X1 U575 ( .A1(n449), .A2(n448), .ZN(n472) );
  BUF_X1 U576 ( .A(n503), .Z(n473) );
  XNOR2_X1 U577 ( .A(n464), .B(n516), .ZN(n450) );
  XNOR2_X1 U578 ( .A(n472), .B(KEYINPUT45), .ZN(n674) );
  BUF_X1 U579 ( .A(n674), .Z(n471) );
  INV_X1 U580 ( .A(n710), .ZN(n452) );
  OR2_X1 U581 ( .A1(n454), .A2(n489), .ZN(n453) );
  INV_X1 U582 ( .A(n488), .ZN(n454) );
  AND2_X1 U583 ( .A1(n493), .A2(n488), .ZN(n455) );
  AND2_X2 U584 ( .A1(n457), .A2(n403), .ZN(n456) );
  AND2_X2 U585 ( .A1(n457), .A2(n403), .ZN(n747) );
  XNOR2_X1 U586 ( .A(n475), .B(n474), .ZN(n643) );
  XOR2_X1 U587 ( .A(n466), .B(G104), .Z(n592) );
  NAND2_X1 U588 ( .A1(n747), .A2(G472), .ZN(n486) );
  NAND2_X1 U589 ( .A1(n747), .A2(G478), .ZN(n512) );
  NAND2_X1 U590 ( .A1(n485), .A2(n462), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n486), .B(n411), .ZN(n485) );
  NAND2_X1 U592 ( .A1(n510), .A2(n462), .ZN(n509) );
  XNOR2_X1 U593 ( .A(n512), .B(n511), .ZN(n510) );
  XNOR2_X1 U594 ( .A(n484), .B(n415), .ZN(G57) );
  XNOR2_X1 U595 ( .A(n459), .B(n458), .ZN(G60) );
  NAND2_X1 U596 ( .A1(n461), .A2(n462), .ZN(n459) );
  XNOR2_X1 U597 ( .A(n460), .B(n414), .ZN(G51) );
  NAND2_X1 U598 ( .A1(n463), .A2(n462), .ZN(n460) );
  NAND2_X1 U599 ( .A1(n621), .A2(n490), .ZN(n488) );
  XNOR2_X1 U600 ( .A(n745), .B(n410), .ZN(n461) );
  XNOR2_X1 U601 ( .A(n738), .B(n412), .ZN(n463) );
  XNOR2_X2 U602 ( .A(n564), .B(n563), .ZN(n752) );
  INV_X4 U603 ( .A(G953), .ZN(n770) );
  XNOR2_X2 U604 ( .A(n623), .B(KEYINPUT105), .ZN(n688) );
  XOR2_X2 U605 ( .A(KEYINPUT10), .B(n536), .Z(n768) );
  XNOR2_X1 U606 ( .A(n538), .B(n519), .ZN(n539) );
  NOR2_X1 U607 ( .A1(n710), .A2(n476), .ZN(n475) );
  XNOR2_X2 U608 ( .A(n545), .B(n546), .ZN(n710) );
  INV_X1 U609 ( .A(KEYINPUT44), .ZN(n490) );
  XOR2_X2 U610 ( .A(KEYINPUT67), .B(G101), .Z(n555) );
  XNOR2_X1 U611 ( .A(n540), .B(n539), .ZN(n749) );
  XNOR2_X2 U612 ( .A(G125), .B(G146), .ZN(n565) );
  NOR2_X2 U613 ( .A1(n615), .A2(n712), .ZN(n627) );
  XNOR2_X2 U614 ( .A(n494), .B(G143), .ZN(n566) );
  NOR2_X2 U615 ( .A1(n503), .A2(n581), .ZN(n582) );
  XNOR2_X2 U616 ( .A(n658), .B(KEYINPUT19), .ZN(n503) );
  XNOR2_X2 U617 ( .A(n506), .B(n504), .ZN(n564) );
  XNOR2_X2 U618 ( .A(n507), .B(n527), .ZN(n506) );
  XNOR2_X2 U619 ( .A(G119), .B(G113), .ZN(n507) );
  XNOR2_X1 U620 ( .A(n509), .B(n508), .ZN(G63) );
  INV_X1 U621 ( .A(n746), .ZN(n511) );
  XNOR2_X2 U622 ( .A(n515), .B(n514), .ZN(n779) );
  NAND2_X1 U623 ( .A1(n613), .A2(n612), .ZN(n515) );
  XNOR2_X1 U624 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n518) );
  AND2_X1 U625 ( .A1(n601), .A2(G221), .ZN(n519) );
  AND2_X1 U626 ( .A1(G210), .A2(n573), .ZN(n520) );
  INV_X1 U627 ( .A(KEYINPUT86), .ZN(n574) );
  NOR2_X1 U628 ( .A1(G952), .A2(n770), .ZN(n521) );
  XOR2_X1 U629 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n530) );
  XOR2_X1 U630 ( .A(n555), .B(KEYINPUT5), .Z(n523) );
  NAND2_X1 U631 ( .A1(n588), .A2(G210), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U633 ( .A(n548), .B(KEYINPUT23), .ZN(n534) );
  XOR2_X1 U634 ( .A(KEYINPUT95), .B(G119), .Z(n532) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U637 ( .A(n535), .B(KEYINPUT24), .Z(n540) );
  XNOR2_X1 U638 ( .A(n768), .B(KEYINPUT73), .ZN(n538) );
  NAND2_X1 U639 ( .A1(G234), .A2(n770), .ZN(n537) );
  XOR2_X1 U640 ( .A(KEYINPUT8), .B(n537), .Z(n601) );
  XOR2_X1 U641 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n543) );
  NAND2_X1 U642 ( .A1(n572), .A2(G234), .ZN(n541) );
  XNOR2_X1 U643 ( .A(n541), .B(KEYINPUT20), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n583), .A2(G217), .ZN(n542) );
  XNOR2_X1 U645 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U646 ( .A(KEYINPUT96), .B(n544), .ZN(n545) );
  NAND2_X1 U647 ( .A1(G227), .A2(n770), .ZN(n550) );
  INV_X1 U648 ( .A(KEYINPUT77), .ZN(n549) );
  INV_X1 U649 ( .A(n552), .ZN(n554) );
  XNOR2_X2 U650 ( .A(n753), .B(n556), .ZN(n567) );
  XNOR2_X1 U651 ( .A(G146), .B(KEYINPUT94), .ZN(n557) );
  XNOR2_X1 U652 ( .A(KEYINPUT71), .B(G469), .ZN(n558) );
  XNOR2_X2 U653 ( .A(n559), .B(n558), .ZN(n645) );
  INV_X1 U654 ( .A(KEYINPUT1), .ZN(n560) );
  XNOR2_X2 U655 ( .A(n645), .B(n560), .ZN(n615) );
  OR2_X1 U656 ( .A1(n615), .A2(n637), .ZN(n561) );
  NOR2_X1 U657 ( .A1(n710), .A2(n561), .ZN(n562) );
  XNOR2_X1 U658 ( .A(KEYINPUT78), .B(n562), .ZN(n612) );
  XNOR2_X1 U659 ( .A(KEYINPUT22), .B(KEYINPUT66), .ZN(n611) );
  NAND2_X1 U660 ( .A1(G224), .A2(n770), .ZN(n568) );
  XNOR2_X1 U661 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U662 ( .A(KEYINPUT4), .B(n570), .ZN(n571) );
  NAND2_X1 U663 ( .A1(G214), .A2(n573), .ZN(n700) );
  NAND2_X1 U664 ( .A1(G237), .A2(G234), .ZN(n575) );
  XNOR2_X1 U665 ( .A(n575), .B(KEYINPUT14), .ZN(n577) );
  NAND2_X1 U666 ( .A1(G952), .A2(n577), .ZN(n576) );
  XOR2_X1 U667 ( .A(KEYINPUT92), .B(n576), .Z(n729) );
  NAND2_X1 U668 ( .A1(n770), .A2(n729), .ZN(n634) );
  NAND2_X1 U669 ( .A1(G902), .A2(n577), .ZN(n632) );
  INV_X1 U670 ( .A(n632), .ZN(n578) );
  NOR2_X1 U671 ( .A1(G898), .A2(n770), .ZN(n756) );
  NAND2_X1 U672 ( .A1(n578), .A2(n756), .ZN(n579) );
  NAND2_X1 U673 ( .A1(n634), .A2(n579), .ZN(n580) );
  XNOR2_X1 U674 ( .A(KEYINPUT93), .B(n580), .ZN(n581) );
  NAND2_X1 U675 ( .A1(n583), .A2(G221), .ZN(n584) );
  XOR2_X1 U676 ( .A(KEYINPUT21), .B(n584), .Z(n709) );
  XNOR2_X1 U677 ( .A(n709), .B(KEYINPUT98), .ZN(n614) );
  XNOR2_X1 U678 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U679 ( .A(n768), .B(n587), .Z(n590) );
  NAND2_X1 U680 ( .A1(n588), .A2(G214), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n590), .B(n589), .ZN(n598) );
  XNOR2_X1 U682 ( .A(n592), .B(n591), .ZN(n596) );
  XNOR2_X1 U683 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n593) );
  XNOR2_X1 U684 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U685 ( .A(n596), .B(n595), .Z(n597) );
  XNOR2_X1 U686 ( .A(n598), .B(n597), .ZN(n744) );
  NOR2_X1 U687 ( .A1(G902), .A2(n744), .ZN(n600) );
  XNOR2_X1 U688 ( .A(KEYINPUT13), .B(G475), .ZN(n599) );
  XNOR2_X1 U689 ( .A(n600), .B(n599), .ZN(n625) );
  NAND2_X1 U690 ( .A1(G217), .A2(n601), .ZN(n602) );
  XNOR2_X1 U691 ( .A(G107), .B(n604), .ZN(n605) );
  XNOR2_X1 U692 ( .A(n606), .B(n605), .ZN(n607) );
  XOR2_X1 U693 ( .A(n608), .B(n607), .Z(n746) );
  NOR2_X1 U694 ( .A1(n746), .A2(G902), .ZN(n609) );
  XOR2_X1 U695 ( .A(G478), .B(n609), .Z(n622) );
  NOR2_X1 U696 ( .A1(n625), .A2(n622), .ZN(n646) );
  XNOR2_X2 U697 ( .A(n616), .B(KEYINPUT33), .ZN(n707) );
  NAND2_X1 U698 ( .A1(n617), .A2(n707), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n625), .A2(n622), .ZN(n663) );
  INV_X1 U700 ( .A(KEYINPUT85), .ZN(n621) );
  INV_X1 U701 ( .A(n622), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n624), .A2(n625), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n691) );
  NOR2_X1 U704 ( .A1(n688), .A2(n691), .ZN(n699) );
  XOR2_X1 U705 ( .A(n699), .B(KEYINPUT81), .Z(n667) );
  INV_X1 U706 ( .A(n712), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n645), .A2(n626), .ZN(n650) );
  NAND2_X1 U708 ( .A1(n715), .A2(n627), .ZN(n720) );
  NAND2_X1 U709 ( .A1(n674), .A2(n354), .ZN(n630) );
  INV_X1 U710 ( .A(n615), .ZN(n640) );
  NOR2_X1 U711 ( .A1(G900), .A2(n632), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G953), .A2(n633), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U714 ( .A(n636), .B(KEYINPUT79), .ZN(n651) );
  NAND2_X1 U715 ( .A1(n688), .A2(n637), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n643), .A2(n638), .ZN(n657) );
  NAND2_X1 U717 ( .A1(n657), .A2(n700), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n641), .B(KEYINPUT43), .ZN(n642) );
  NOR2_X1 U720 ( .A1(n501), .A2(n642), .ZN(n696) );
  XOR2_X1 U721 ( .A(KEYINPUT38), .B(n501), .Z(n701) );
  NAND2_X1 U722 ( .A1(n701), .A2(n700), .ZN(n698) );
  INV_X1 U723 ( .A(n646), .ZN(n703) );
  NOR2_X1 U724 ( .A1(n698), .A2(n703), .ZN(n647) );
  XOR2_X1 U725 ( .A(KEYINPUT41), .B(n647), .Z(n723) );
  NAND2_X1 U726 ( .A1(n666), .A2(n723), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT42), .ZN(n783) );
  INV_X1 U728 ( .A(n701), .ZN(n653) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U730 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n672) );
  NAND2_X1 U732 ( .A1(n688), .A2(n672), .ZN(n656) );
  AND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT36), .B(n659), .Z(n660) );
  NOR2_X1 U735 ( .A1(n615), .A2(n660), .ZN(n693) );
  INV_X1 U736 ( .A(n631), .ZN(n662) );
  NAND2_X1 U737 ( .A1(KEYINPUT47), .A2(n699), .ZN(n664) );
  XOR2_X1 U738 ( .A(KEYINPUT80), .B(n664), .Z(n665) );
  NOR2_X1 U739 ( .A1(n781), .A2(n665), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n686), .A2(n667), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n691), .ZN(n695) );
  NAND2_X1 U743 ( .A1(n354), .A2(KEYINPUT2), .ZN(n673) );
  INV_X1 U744 ( .A(KEYINPUT2), .ZN(n675) );
  XOR2_X1 U745 ( .A(G104), .B(KEYINPUT111), .Z(n677) );
  NAND2_X1 U746 ( .A1(n678), .A2(n688), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n677), .B(n676), .ZN(G6) );
  XOR2_X1 U748 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n680) );
  NAND2_X1 U749 ( .A1(n678), .A2(n691), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U751 ( .A(G107), .B(n681), .ZN(G9) );
  XOR2_X1 U752 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n683) );
  NAND2_X1 U753 ( .A1(n691), .A2(n686), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n685) );
  XOR2_X1 U755 ( .A(G128), .B(KEYINPUT112), .Z(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(G30) );
  NAND2_X1 U757 ( .A1(n686), .A2(n688), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(G146), .ZN(G48) );
  XOR2_X1 U759 ( .A(n466), .B(KEYINPUT115), .Z(n690) );
  XNOR2_X1 U760 ( .A(n690), .B(n689), .ZN(G15) );
  XNOR2_X1 U761 ( .A(n692), .B(G116), .ZN(G18) );
  XNOR2_X1 U762 ( .A(G125), .B(n693), .ZN(n694) );
  XNOR2_X1 U763 ( .A(n694), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U764 ( .A(G134), .B(n695), .ZN(G36) );
  XOR2_X1 U765 ( .A(G140), .B(n696), .Z(G42) );
  XOR2_X1 U766 ( .A(KEYINPUT2), .B(n697), .Z(n735) );
  NAND2_X1 U767 ( .A1(n723), .A2(n707), .ZN(n732) );
  OR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n706) );
  NOR2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT118), .B(n704), .Z(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n726) );
  NOR2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U775 ( .A(KEYINPUT49), .B(n711), .ZN(n718) );
  XOR2_X1 U776 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n714) );
  NAND2_X1 U777 ( .A1(n615), .A2(n712), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n721), .B(KEYINPUT51), .ZN(n722) );
  XNOR2_X1 U783 ( .A(n722), .B(KEYINPUT117), .ZN(n724) );
  NAND2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n728) );
  XOR2_X1 U786 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n727) );
  XNOR2_X1 U787 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U788 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U789 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U790 ( .A(KEYINPUT120), .B(n733), .Z(n734) );
  NAND2_X1 U791 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U792 ( .A1(n736), .A2(G953), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n737), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U794 ( .A1(n747), .A2(G210), .ZN(n738) );
  XOR2_X1 U795 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n740) );
  NAND2_X1 U796 ( .A1(n402), .A2(G469), .ZN(n739) );
  NOR2_X1 U797 ( .A1(n751), .A2(n742), .ZN(G54) );
  NAND2_X1 U798 ( .A1(n456), .A2(G475), .ZN(n745) );
  INV_X1 U799 ( .A(KEYINPUT59), .ZN(n743) );
  NAND2_X1 U800 ( .A1(G217), .A2(n402), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n751), .A2(n750), .ZN(G66) );
  BUF_X1 U803 ( .A(n752), .Z(n755) );
  XOR2_X1 U804 ( .A(n753), .B(G101), .Z(n754) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(n757) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n766) );
  XOR2_X1 U807 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n759) );
  NAND2_X1 U808 ( .A1(G224), .A2(G953), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U810 ( .A1(G898), .A2(n760), .ZN(n761) );
  XNOR2_X1 U811 ( .A(n761), .B(KEYINPUT124), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n471), .A2(n770), .ZN(n762) );
  NAND2_X1 U813 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U814 ( .A(n764), .B(KEYINPUT125), .Z(n765) );
  XNOR2_X1 U815 ( .A(n766), .B(n765), .ZN(G69) );
  XNOR2_X1 U816 ( .A(n768), .B(n767), .ZN(n772) );
  INV_X1 U817 ( .A(n772), .ZN(n769) );
  NAND2_X1 U818 ( .A1(n771), .A2(n770), .ZN(n777) );
  XOR2_X1 U819 ( .A(n772), .B(G227), .Z(n773) );
  XNOR2_X1 U820 ( .A(n773), .B(KEYINPUT126), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U822 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U824 ( .A(n778), .B(G122), .Z(G24) );
  XNOR2_X1 U825 ( .A(G119), .B(KEYINPUT127), .ZN(n780) );
  XNOR2_X1 U826 ( .A(n780), .B(n779), .ZN(G21) );
  XOR2_X1 U827 ( .A(G143), .B(n781), .Z(n782) );
  XNOR2_X1 U828 ( .A(KEYINPUT114), .B(n782), .ZN(G45) );
  XNOR2_X1 U829 ( .A(G137), .B(n783), .ZN(G39) );
endmodule

