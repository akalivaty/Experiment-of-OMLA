//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n437, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1238, new_n1239,
    new_n1240, new_n1241;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  INV_X1    g010(.A(G132), .ZN(G219));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G82), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n434), .A2(new_n437), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G136), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n481), .A2(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(G114), .B2(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n494), .B(new_n496), .C1(new_n469), .C2(new_n468), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n468), .B2(new_n469), .ZN(new_n498));
  INV_X1    g073(.A(new_n496), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n492), .B1(new_n497), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n506), .A2(new_n509), .A3(G88), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n510), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT7), .Z(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(G51), .B2(new_n511), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n506), .A2(new_n509), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n506), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n504), .A2(KEYINPUT72), .A3(new_n505), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n527), .A2(G64), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n514), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  NAND3_X1  g111(.A1(new_n524), .A2(G56), .A3(new_n525), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n514), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n511), .A2(G43), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n521), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT75), .Z(G188));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n504), .B2(new_n505), .ZN(new_n552));
  AND2_X1   g127(.A1(G78), .A2(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT78), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n556), .B(G651), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  INV_X1    g132(.A(new_n521), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n555), .A2(new_n557), .B1(G91), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n511), .A2(G53), .ZN(new_n561));
  AND2_X1   g136(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n562));
  NOR2_X1   g137(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n511), .B2(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n566), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n511), .B(G53), .C1(new_n562), .C2(new_n563), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(KEYINPUT77), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n559), .A2(new_n567), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n514), .B1(new_n526), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n511), .A2(G49), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n521), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n511), .A2(G48), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n521), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n506), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n514), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n526), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n511), .A2(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n521), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n592), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(new_n506), .A2(G66), .ZN(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n503), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n601));
  NAND3_X1  g176(.A1(new_n558), .A2(G92), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n601), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n521), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n600), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G321));
  NOR2_X1   g185(.A1(G168), .A2(new_n607), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n607), .B2(G299), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(G297));
  XOR2_X1   g188(.A(new_n612), .B(KEYINPUT81), .Z(G280));
  INV_X1    g189(.A(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  INV_X1    g192(.A(new_n543), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n607), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n606), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n464), .A2(new_n472), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT13), .Z(new_n625));
  XOR2_X1   g200(.A(KEYINPUT82), .B(G2100), .Z(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT83), .Z(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n478), .A2(G123), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT84), .ZN(new_n633));
  AOI211_X1 g208(.A(new_n631), .B(new_n633), .C1(G135), .C2(new_n485), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n626), .A2(new_n625), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n628), .B(new_n636), .C1(new_n635), .C2(new_n634), .ZN(G156));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n638), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(KEYINPUT86), .A3(KEYINPUT14), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n644), .A2(new_n645), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n642), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI211_X1 g229(.A(new_n652), .B(new_n641), .C1(new_n649), .C2(new_n650), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n640), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n650), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT86), .B1(new_n646), .B2(KEYINPUT14), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(new_n641), .ZN(new_n660));
  INV_X1    g235(.A(new_n640), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n651), .A2(new_n653), .A3(new_n642), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(new_n656), .B2(new_n663), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  NOR3_X1   g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n702), .ZN(new_n705));
  INV_X1    g280(.A(new_n699), .ZN(new_n706));
  INV_X1    g281(.A(new_n698), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n696), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n705), .B1(new_n708), .B2(new_n700), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G22), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n712), .A2(G6), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n587), .B2(new_n712), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT32), .B(G1981), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n712), .A2(G23), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n579), .B2(new_n712), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT33), .B(G1976), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n715), .A2(G24), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n592), .A2(new_n595), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n715), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1986), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G25), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT89), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n485), .A2(G131), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n478), .A2(G119), .ZN(new_n742));
  OR2_X1    g317(.A1(G95), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n732), .A2(new_n733), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT36), .ZN(new_n751));
  NOR2_X1   g326(.A1(G162), .A2(new_n738), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n738), .B2(G35), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n755), .A2(KEYINPUT98), .A3(G2090), .ZN(new_n756));
  INV_X1    g331(.A(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n464), .A2(G2105), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n464), .A2(new_n463), .ZN(new_n759));
  INV_X1    g334(.A(G140), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n471), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n738), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n738), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n712), .A2(G4), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n615), .B2(new_n712), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1348), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n738), .A2(G32), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G129), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT26), .Z(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT97), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n782), .A2(new_n788), .A3(new_n783), .A4(new_n785), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n781), .B1(new_n791), .B2(new_n738), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT27), .B(G1996), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n780), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n715), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G20), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT23), .ZN(new_n798));
  INV_X1    g373(.A(G299), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n712), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT100), .B(G1956), .Z(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n756), .A2(new_n777), .A3(new_n795), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n738), .A2(G33), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT25), .Z(new_n806));
  INV_X1    g381(.A(G139), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n759), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n463), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n804), .B1(new_n811), .B2(new_n738), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G2072), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT96), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(G2072), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G11), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(G11), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(G28), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n738), .B1(new_n819), .B2(G28), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n817), .B(new_n818), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n634), .B2(G29), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT24), .ZN(new_n824));
  INV_X1    g399(.A(G34), .ZN(new_n825));
  AOI21_X1  g400(.A(G29), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G160), .B2(new_n738), .ZN(new_n828));
  INV_X1    g403(.A(G2084), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n814), .A2(new_n815), .A3(new_n823), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n712), .A2(G21), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G168), .B2(new_n712), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(G1966), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(G1966), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n738), .A2(G27), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G164), .B2(new_n738), .ZN(new_n837));
  INV_X1    g412(.A(G2078), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n712), .A2(G5), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G171), .B2(new_n712), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1961), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n831), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n753), .B(KEYINPUT29), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n846));
  INV_X1    g421(.A(G2090), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT99), .B1(new_n755), .B2(G2090), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT98), .B1(new_n755), .B2(G2090), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n800), .A2(new_n801), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n796), .A2(G19), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT92), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n543), .B2(new_n796), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(G1341), .Z(new_n856));
  NAND3_X1  g431(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n803), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n751), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(G311));
  XNOR2_X1  g435(.A(new_n859), .B(KEYINPUT101), .ZN(G150));
  NAND2_X1  g436(.A1(new_n615), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n524), .A2(G67), .A3(new_n525), .ZN(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n514), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n511), .A2(G55), .ZN(new_n867));
  INV_X1    g442(.A(G93), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n521), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n618), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n543), .A2(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n863), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n876));
  AOI21_X1  g451(.A(G860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(G860), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT37), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT102), .ZN(G145));
  NAND2_X1  g457(.A1(new_n481), .A2(new_n486), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G160), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n634), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT106), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n478), .A2(G130), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n463), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(G142), .B2(new_n485), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(new_n624), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n745), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n770), .B1(new_n787), .B2(new_n789), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n811), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n770), .A2(new_n787), .A3(new_n789), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n811), .B1(new_n899), .B2(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G114), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n489), .B1(new_n902), .B2(G2105), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(G126), .B2(new_n478), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n500), .A2(new_n905), .A3(new_n497), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n500), .B2(new_n497), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n497), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n496), .B1(new_n464), .B2(new_n494), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT103), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n500), .A2(new_n905), .A3(new_n497), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n492), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n898), .A2(new_n900), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n886), .B1(new_n893), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  INV_X1    g493(.A(new_n915), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n914), .B1(new_n898), .B2(new_n900), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n909), .A2(new_n922), .A3(new_n915), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n893), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g501(.A(KEYINPUT105), .B(new_n893), .C1(new_n921), .C2(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n917), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n916), .B(new_n893), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n929), .B2(new_n885), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n874), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n620), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G299), .A2(new_n606), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G299), .A2(new_n606), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n938), .B2(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n934), .B(new_n620), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(new_n940), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT42), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G290), .A2(new_n587), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n735), .A2(G305), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G288), .A2(G166), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n579), .A2(G303), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n951), .A2(new_n954), .A3(new_n955), .A4(new_n952), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n948), .A2(new_n945), .A3(new_n942), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n950), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n950), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n871), .A2(new_n607), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(G295));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n968), .ZN(G331));
  NAND2_X1  g545(.A1(new_n874), .A2(G171), .ZN(new_n971));
  NAND3_X1  g546(.A1(G301), .A2(new_n872), .A3(new_n873), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(G168), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G168), .B1(new_n971), .B2(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n940), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G286), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n946), .A2(new_n978), .A3(new_n973), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n979), .A3(new_n959), .ZN(new_n980));
  INV_X1    g555(.A(G37), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n959), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n957), .A2(KEYINPUT110), .A3(new_n958), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n979), .B2(new_n976), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n986), .ZN(new_n989));
  INV_X1    g564(.A(new_n939), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n937), .A3(new_n943), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n991), .A2(KEYINPUT111), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT41), .B1(new_n938), .B2(new_n939), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n991), .A3(KEYINPUT111), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n992), .A2(new_n978), .A3(new_n973), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n976), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n981), .A4(new_n980), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n988), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n982), .ZN(new_n1003));
  INV_X1    g578(.A(new_n987), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT43), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n986), .B1(new_n976), .B2(new_n995), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n982), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n997), .A2(KEYINPUT112), .A3(new_n981), .A4(new_n980), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1005), .B1(new_n1010), .B2(KEYINPUT43), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1002), .B1(new_n1011), .B2(new_n1001), .ZN(G397));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n908), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n467), .A2(new_n1015), .A3(new_n474), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n770), .B(G2067), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n790), .A2(G1996), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n790), .A2(G1996), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n747), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n745), .B(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1018), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G290), .B(G1986), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1018), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT113), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(G1384), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1016), .B1(G164), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n908), .A2(new_n1013), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n1030), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n1035), .B2(G1966), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n500), .A2(new_n497), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n1037), .B2(new_n904), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1016), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n914), .A2(G1384), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1039), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n829), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1044), .B(new_n1045), .C1(new_n1014), .C2(new_n1033), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1036), .A2(G168), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1033), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1030), .B1(new_n914), .B2(G1384), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1966), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1051), .A2(new_n1044), .B1(new_n1042), .B2(new_n829), .ZN(new_n1052));
  AOI21_X1  g627(.A(G168), .B1(new_n1052), .B2(new_n1036), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT51), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1047), .A2(new_n1056), .A3(G8), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  INV_X1    g637(.A(new_n474), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n465), .A2(new_n466), .ZN(new_n1064));
  OAI211_X1 g639(.A(G40), .B(new_n1063), .C1(new_n1064), .C2(new_n463), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1037), .A2(new_n904), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1013), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(new_n1067), .B2(KEYINPUT50), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n847), .C1(new_n1034), .C2(KEYINPUT50), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n914), .A2(new_n1032), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1016), .B1(new_n1038), .B2(KEYINPUT45), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT114), .B(new_n718), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g648(.A(new_n1016), .B1(new_n1038), .B2(KEYINPUT45), .C1(new_n914), .C2(new_n1032), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT114), .B1(new_n1074), .B2(new_n718), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1062), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G303), .A2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT116), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  NAND4_X1  g655(.A1(G303), .A2(new_n1080), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT117), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1077), .A2(KEYINPUT117), .A3(new_n1078), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n718), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT115), .A3(new_n1072), .A4(new_n1069), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1076), .A2(G8), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT50), .B1(new_n914), .B2(G1384), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1065), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n847), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1086), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1085), .B1(new_n1094), .B2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(G1976), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(G288), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n908), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n579), .A2(G1976), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1097), .A2(G8), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n587), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(G1981), .B1(new_n583), .B2(new_n586), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT49), .A3(new_n1103), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(G8), .A3(new_n1098), .A4(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1098), .A2(new_n1099), .A3(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT52), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1100), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1095), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1068), .B1(new_n1034), .B2(KEYINPUT50), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1961), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1068), .B(KEYINPUT121), .C1(new_n1034), .C2(KEYINPUT50), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1035), .A2(KEYINPUT53), .A3(new_n838), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1074), .B2(G2078), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1090), .A2(new_n1112), .A3(G171), .A4(new_n1122), .ZN(new_n1123));
  NOR4_X1   g698(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(KEYINPUT62), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT125), .B1(new_n1126), .B2(new_n1058), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1076), .A2(G8), .A3(new_n1089), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1085), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G168), .A2(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1052), .B2(new_n1036), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1111), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1090), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1090), .A2(new_n1112), .A3(new_n1133), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(KEYINPUT120), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1134), .B1(new_n1137), .B2(KEYINPUT120), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1108), .A2(new_n1141), .B1(new_n1101), .B2(new_n587), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  OAI211_X1 g718(.A(G8), .B(new_n1098), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1090), .A2(new_n1111), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(G1956), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1039), .B1(new_n908), .B2(new_n1013), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1016), .B1(new_n1067), .B2(KEYINPUT50), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n568), .B2(new_n569), .ZN(new_n1152));
  AOI22_X1  g727(.A1(G299), .A2(KEYINPUT57), .B1(new_n559), .B2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT56), .B(G2072), .Z(new_n1154));
  OAI211_X1 g729(.A(new_n1151), .B(new_n1153), .C1(new_n1074), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G1348), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1115), .A2(new_n1157), .A3(new_n1117), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1041), .A2(new_n776), .A3(new_n1016), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n615), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n559), .A2(new_n1152), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(G1956), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1070), .A2(new_n1071), .A3(new_n1154), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1156), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1070), .A2(new_n1071), .A3(G1996), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT58), .B(G1341), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1041), .B2(new_n1016), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n543), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1174), .B(new_n543), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1167), .A2(new_n1155), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1167), .B2(new_n1155), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1160), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n615), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1158), .A2(KEYINPUT60), .A3(new_n1159), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT122), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1158), .A2(new_n1186), .A3(KEYINPUT60), .A4(new_n1159), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1180), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1185), .A2(new_n1182), .A3(new_n615), .A4(new_n1187), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1168), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1122), .A2(G171), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1063), .A2(KEYINPUT123), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1193), .A2(new_n1015), .A3(new_n467), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n474), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1196), .A2(new_n1014), .A3(KEYINPUT124), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT124), .B1(new_n1196), .B2(new_n1014), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1070), .A2(new_n1120), .A3(G2078), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1118), .B(new_n1121), .C1(new_n1197), .C2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1192), .B1(G171), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT54), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1201), .A2(G171), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1205), .B(KEYINPUT54), .C1(G171), .C2(new_n1122), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1090), .A2(new_n1112), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1204), .A2(new_n1206), .A3(new_n1125), .A4(new_n1207), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1140), .B(new_n1147), .C1(new_n1191), .C2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1029), .B1(new_n1128), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(G290), .A2(G1986), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT48), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1212), .A2(new_n1213), .A3(new_n1017), .ZN(new_n1214));
  AOI21_X1  g789(.A(KEYINPUT48), .B1(new_n1211), .B2(new_n1018), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1026), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1017), .A2(G1996), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT46), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1017), .B1(new_n1019), .B2(new_n791), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT47), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n770), .A2(new_n776), .ZN(new_n1222));
  OR2_X1    g797(.A1(new_n745), .A2(new_n1023), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1022), .B2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g799(.A(new_n1216), .B(new_n1221), .C1(new_n1018), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1210), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g801(.A1(new_n461), .A2(G227), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n666), .B2(new_n667), .ZN(new_n1229));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g805(.A(new_n1228), .B(KEYINPUT126), .C1(new_n666), .C2(new_n667), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1231), .A2(new_n710), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g807(.A(new_n1233), .B1(new_n928), .B2(new_n930), .ZN(new_n1234));
  AND3_X1   g808(.A1(new_n1000), .A2(new_n1234), .A3(KEYINPUT127), .ZN(new_n1235));
  AOI21_X1  g809(.A(KEYINPUT127), .B1(new_n1000), .B2(new_n1234), .ZN(new_n1236));
  NOR2_X1   g810(.A1(new_n1235), .A2(new_n1236), .ZN(G308));
  NAND2_X1  g811(.A1(new_n1000), .A2(new_n1234), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n1234), .A3(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1241), .ZN(G225));
endmodule


