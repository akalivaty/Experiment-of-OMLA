//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  AOI21_X1  g000(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G127gat), .A2(G134gat), .ZN(new_n206));
  OAI221_X1 g005(.A(new_n202), .B1(G113gat), .B2(G120gat), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n202), .B1(G113gat), .B2(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n206), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT70), .B(G134gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n203), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n208), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT27), .B(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n217), .A2(new_n218), .B1(new_n219), .B2(KEYINPUT28), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n220), .A2(new_n219), .A3(KEYINPUT28), .ZN(new_n221));
  AND2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT26), .ZN(new_n226));
  AOI211_X1 g025(.A(new_n222), .B(new_n226), .C1(KEYINPUT26), .C2(new_n225), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n220), .B1(new_n219), .B2(KEYINPUT28), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n225), .B2(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n224), .B1(KEYINPUT23), .B2(new_n225), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(KEYINPUT67), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT23), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n223), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n239), .B2(new_n240), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n236), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT67), .B1(new_n243), .B2(new_n245), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n231), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n243), .A2(new_n245), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n246), .A4(new_n252), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n230), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n216), .B1(new_n260), .B2(KEYINPUT72), .ZN(new_n261));
  AND4_X1   g060(.A1(KEYINPUT25), .A2(new_n236), .A3(new_n241), .A4(new_n242), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n244), .B1(new_n251), .B2(new_n236), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(KEYINPUT67), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT68), .B1(new_n264), .B2(new_n258), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n253), .A2(new_n231), .A3(new_n254), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n229), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT64), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n216), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT32), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT33), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G15gat), .B(G43gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT73), .ZN(new_n279));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  AOI21_X1  g080(.A(new_n275), .B1(new_n281), .B2(KEYINPUT33), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n277), .A2(new_n281), .B1(new_n274), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT34), .ZN(new_n284));
  INV_X1    g083(.A(new_n272), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(KEYINPUT75), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n273), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n285), .ZN(new_n289));
  AOI211_X1 g088(.A(new_n272), .B(new_n286), .C1(new_n270), .C2(new_n273), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G155gat), .B(G162gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT80), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT79), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(G141gat), .ZN(new_n298));
  INV_X1    g097(.A(G141gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n300), .C1(new_n299), .C2(G148gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G155gat), .B(G162gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT2), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n295), .A2(new_n301), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n294), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(KEYINPUT22), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G211gat), .B(G218gat), .Z(new_n318));
  AND2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n317), .A2(new_n318), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n312), .B1(new_n322), .B2(KEYINPUT3), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G228gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G22gat), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n323), .A2(new_n325), .A3(G228gat), .A4(G233gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT31), .B(G50gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT84), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n329), .A2(new_n331), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n340), .A2(new_n330), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT84), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n334), .A2(new_n342), .A3(new_n337), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n339), .A2(new_n332), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n332), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n334), .B2(new_n337), .ZN(new_n346));
  INV_X1    g145(.A(new_n337), .ZN(new_n347));
  AOI211_X1 g146(.A(KEYINPUT84), .B(new_n347), .C1(new_n332), .C2(new_n333), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n283), .A2(new_n291), .A3(KEYINPUT76), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT76), .B1(new_n283), .B2(new_n291), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n293), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G226gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n328), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT29), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n229), .B1(new_n254), .B2(new_n253), .ZN(new_n362));
  INV_X1    g161(.A(new_n359), .ZN(new_n363));
  OAI22_X1  g162(.A1(new_n260), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n321), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n360), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n267), .B2(new_n363), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n368), .B2(new_n365), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n357), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(new_n370), .A3(new_n366), .A4(new_n356), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT30), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n366), .A2(new_n370), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n374), .A4(new_n356), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n214), .A2(new_n215), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n207), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  INV_X1    g185(.A(new_n312), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n216), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n383), .A2(new_n312), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT5), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT81), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n391), .B1(new_n383), .B2(new_n312), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n385), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n216), .A2(new_n387), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n390), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(KEYINPUT5), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n398), .A2(new_n404), .A3(new_n409), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT35), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n353), .A2(new_n380), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n277), .A2(new_n281), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n274), .A2(new_n282), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(KEYINPUT74), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT74), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n274), .A2(new_n282), .ZN(new_n424));
  INV_X1    g223(.A(new_n281), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n274), .B2(new_n276), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n289), .A2(new_n290), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n376), .A2(new_n379), .B1(new_n414), .B2(new_n415), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT35), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n283), .A2(new_n291), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n283), .A2(new_n291), .A3(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(new_n429), .A3(new_n431), .A4(new_n350), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n419), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n431), .A2(new_n350), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n374), .A2(new_n445), .A3(new_n370), .A4(new_n366), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n357), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n377), .B2(new_n374), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT38), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n414), .A2(new_n375), .A3(new_n415), .ZN(new_n452));
  INV_X1    g251(.A(new_n447), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n445), .B1(new_n368), .B2(new_n321), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n364), .A2(new_n321), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT38), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n447), .C2(new_n448), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  OR3_X1    g259(.A1(new_n393), .A2(KEYINPUT39), .A3(new_n397), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n409), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n393), .A2(new_n397), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n390), .A2(new_n402), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT39), .B1(new_n464), .B2(new_n396), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n460), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n411), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n462), .A2(new_n460), .A3(new_n466), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n380), .A2(new_n470), .B1(new_n344), .B2(new_n349), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n444), .B1(new_n459), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n292), .B1(new_n438), .B2(new_n439), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n429), .B1(new_n351), .B2(new_n352), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT36), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n443), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(G57gat), .A2(G64gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(G57gat), .A2(G64gat), .ZN(new_n482));
  AND2_X1   g281(.A1(G71gat), .A2(G78gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(KEYINPUT9), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(KEYINPUT91), .B2(new_n483), .ZN(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G78gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT21), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G231gat), .A2(G233gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G127gat), .B(G155gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT20), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n491), .B(new_n493), .Z(new_n494));
  XOR2_X1   g293(.A(G183gat), .B(G211gat), .Z(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n496), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(G15gat), .B(G22gat), .Z(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT88), .ZN(new_n501));
  INV_X1    g300(.A(G1gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n502), .A2(KEYINPUT16), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n501), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n488), .B2(new_n487), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n499), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT87), .B(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  OR3_X1    g313(.A1(new_n514), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n513), .A2(KEYINPUT15), .A3(new_n515), .A4(new_n516), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT93), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G99gat), .B(G106gat), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(G85gat), .ZN(new_n536));
  INV_X1    g335(.A(G92gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT94), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n538), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n532), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT95), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(KEYINPUT95), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n524), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n546), .ZN(new_n550));
  XOR2_X1   g349(.A(G190gat), .B(G218gat), .Z(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G134gat), .B(G162gat), .Z(new_n555));
  AOI21_X1  g354(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT96), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(KEYINPUT96), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n511), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n539), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n487), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n546), .A2(new_n487), .B1(new_n566), .B2(new_n543), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n546), .A2(new_n568), .A3(new_n487), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  OAI211_X1 g376(.A(new_n574), .B(new_n577), .C1(new_n573), .C2(new_n567), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n567), .A2(new_n573), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n570), .B1(new_n568), .B2(new_n567), .ZN(new_n581));
  INV_X1    g380(.A(new_n573), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n546), .A2(new_n487), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n543), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n584), .A2(new_n568), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(KEYINPUT97), .B(new_n573), .C1(new_n586), .C2(new_n570), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n578), .B1(new_n588), .B2(new_n577), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n564), .A2(KEYINPUT98), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n528), .A2(new_n592), .A3(new_n507), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n507), .A2(new_n549), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G229gat), .A2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n527), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n507), .B1(new_n525), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT89), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n595), .A2(KEYINPUT18), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n596), .A3(new_n593), .A4(new_n594), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT18), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n507), .B(new_n549), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n596), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G197gat), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT11), .B(G169gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n600), .A2(new_n603), .A3(new_n615), .A4(new_n607), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n563), .B2(new_n589), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n591), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n480), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n416), .B(KEYINPUT99), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G1gat), .ZN(G1324gat));
  INV_X1    g423(.A(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n376), .A2(new_n379), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT16), .B(G8gat), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n506), .B1(new_n621), .B2(new_n380), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT42), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(KEYINPUT42), .B2(new_n628), .ZN(G1325gat));
  INV_X1    g430(.A(new_n473), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n625), .A2(G15gat), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n474), .B1(new_n440), .B2(new_n429), .ZN(new_n634));
  AOI211_X1 g433(.A(KEYINPUT36), .B(new_n292), .C1(new_n438), .C2(new_n439), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT100), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n475), .A2(new_n477), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT101), .B1(new_n636), .B2(new_n638), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G15gat), .B1(new_n625), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n633), .A2(new_n645), .ZN(G1326gat));
  INV_X1    g445(.A(new_n350), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n621), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT102), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  INV_X1    g450(.A(new_n562), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n614), .A2(new_n616), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n653), .A2(new_n511), .A3(new_n589), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n652), .B(new_n654), .C1(new_n443), .C2(new_n478), .ZN(new_n655));
  INV_X1    g454(.A(new_n622), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n655), .A2(G29gat), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT45), .Z(new_n658));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n652), .C1(new_n443), .C2(new_n478), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n654), .B(KEYINPUT103), .ZN(new_n660));
  INV_X1    g459(.A(new_n419), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n441), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT86), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n636), .A2(new_n472), .A3(new_n638), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n562), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n659), .B(new_n660), .C1(new_n666), .C2(KEYINPUT44), .ZN(new_n667));
  OAI21_X1  g466(.A(G29gat), .B1(new_n667), .B2(new_n656), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n658), .A2(new_n668), .ZN(G1328gat));
  NOR3_X1   g468(.A1(new_n655), .A2(new_n626), .A3(new_n512), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT46), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n512), .B1(new_n667), .B2(new_n626), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1329gat));
  INV_X1    g472(.A(new_n639), .ZN(new_n674));
  OAI21_X1  g473(.A(G43gat), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n655), .A2(G43gat), .A3(new_n632), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT47), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n667), .A2(new_n644), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n676), .B1(new_n680), .B2(G43gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n681), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g481(.A1(new_n350), .A2(G50gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT48), .B1(new_n655), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n636), .A2(new_n472), .A3(new_n638), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n652), .B1(new_n686), .B2(new_n443), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(new_n647), .A3(new_n659), .A4(new_n660), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT105), .B(new_n685), .C1(new_n690), .C2(G50gat), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  OAI21_X1  g491(.A(G50gat), .B1(new_n667), .B2(new_n350), .ZN(new_n693));
  INV_X1    g492(.A(new_n685), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(G50gat), .C1(new_n667), .C2(new_n350), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT104), .B1(new_n655), .B2(new_n684), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n690), .B2(G50gat), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n691), .A2(new_n695), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI221_X1 g503(.A(KEYINPUT106), .B1(new_n699), .B2(new_n701), .C1(new_n691), .C2(new_n695), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1331gat));
  NAND3_X1  g505(.A1(new_n564), .A2(new_n653), .A3(new_n589), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n664), .B2(new_n665), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n622), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT107), .B(G57gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  AND2_X1   g510(.A1(new_n708), .A2(new_n380), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  AND2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n712), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT108), .ZN(G1333gat));
  NAND3_X1  g516(.A1(new_n643), .A2(G71gat), .A3(new_n708), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n708), .A2(new_n473), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(G71gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g520(.A1(new_n708), .A2(new_n647), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n511), .A2(new_n617), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n689), .A2(new_n589), .A3(new_n659), .A4(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n656), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n666), .A2(new_n724), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT51), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n666), .A2(new_n729), .A3(new_n724), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n730), .A3(new_n589), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n622), .A2(new_n536), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  OAI21_X1  g532(.A(G92gat), .B1(new_n725), .B2(new_n626), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n626), .A2(G92gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n728), .A2(new_n730), .A3(new_n589), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n737), .B2(KEYINPUT110), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n734), .A2(new_n739), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT52), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT109), .B(KEYINPUT52), .C1(new_n737), .C2(KEYINPUT110), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n725), .B2(new_n644), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n632), .A2(G99gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n731), .B2(new_n746), .ZN(G1338gat));
  OR3_X1    g546(.A1(new_n731), .A2(G106gat), .A3(new_n350), .ZN(new_n748));
  OAI21_X1  g547(.A(G106gat), .B1(new_n725), .B2(new_n350), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1339gat));
  INV_X1    g553(.A(new_n511), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n583), .A2(new_n756), .A3(new_n587), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n581), .A2(new_n582), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n574), .A2(new_n758), .A3(KEYINPUT54), .ZN(new_n759));
  INV_X1    g558(.A(new_n577), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n757), .A2(KEYINPUT55), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n578), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n756), .B1(new_n572), .B2(new_n573), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n577), .B1(new_n763), .B2(new_n758), .ZN(new_n764));
  AOI211_X1 g563(.A(KEYINPUT111), .B(KEYINPUT55), .C1(new_n764), .C2(new_n757), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n757), .A2(new_n760), .A3(new_n759), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n617), .B(new_n762), .C1(new_n765), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n596), .B1(new_n595), .B2(new_n599), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n604), .A2(new_n606), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n612), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n616), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n590), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n652), .B1(new_n770), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n578), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n583), .A2(new_n756), .A3(new_n587), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT54), .B1(new_n581), .B2(new_n582), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n586), .A2(new_n573), .A3(new_n570), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n760), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n768), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT111), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n766), .A3(new_n768), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n778), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n562), .A2(new_n774), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n755), .B1(new_n777), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n563), .A2(new_n617), .A3(new_n589), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n656), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n380), .A3(new_n353), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795), .B2(new_n653), .ZN(new_n796));
  INV_X1    g595(.A(new_n430), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT112), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n797), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n380), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT113), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n653), .A2(G113gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n795), .B2(new_n590), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n590), .A2(G120gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n802), .B2(new_n806), .ZN(G1341gat));
  NAND3_X1  g606(.A1(new_n801), .A2(new_n203), .A3(new_n511), .ZN(new_n808));
  OAI21_X1  g607(.A(G127gat), .B1(new_n795), .B2(new_n755), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1342gat));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n652), .A2(new_n211), .ZN(new_n812));
  INV_X1    g611(.A(new_n800), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n626), .B(new_n812), .C1(new_n813), .C2(new_n798), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n814), .B2(KEYINPUT56), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .A3(new_n816), .A4(new_n812), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n204), .B1(new_n794), .B2(new_n652), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n814), .B2(KEYINPUT56), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(KEYINPUT115), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1343gat));
  NOR3_X1   g624(.A1(new_n639), .A2(new_n380), .A3(new_n656), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n647), .A2(KEYINPUT57), .ZN(new_n827));
  INV_X1    g626(.A(new_n788), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n783), .A2(KEYINPUT116), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n767), .A2(new_n830), .A3(new_n768), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n762), .A2(new_n829), .A3(new_n617), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n652), .B1(new_n832), .B2(new_n776), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n755), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n827), .B1(new_n838), .B2(new_n791), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n350), .B1(new_n789), .B2(new_n791), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(KEYINPUT57), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n826), .B(new_n617), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(G141gat), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n643), .B2(new_n350), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n647), .C1(new_n641), .C2(new_n642), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n793), .A2(new_n380), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n653), .A2(G141gat), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT58), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(KEYINPUT58), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n842), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n653), .A2(new_n778), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n829), .A2(new_n831), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n775), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n857), .B2(new_n652), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n836), .A3(new_n828), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n790), .B1(new_n859), .B2(new_n755), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n860), .A2(new_n827), .B1(KEYINPUT57), .B2(new_n840), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n861), .A2(KEYINPUT119), .A3(new_n617), .A4(new_n826), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n862), .A3(G141gat), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n852), .A2(new_n863), .A3(KEYINPUT120), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT120), .B1(new_n852), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(G1344gat));
  AND3_X1   g665(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n297), .A3(new_n589), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n755), .B1(new_n833), .B2(new_n788), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n591), .A2(new_n653), .A3(new_n619), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n870), .B(new_n871), .C1(new_n874), .C2(new_n350), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n840), .A2(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n350), .B1(new_n872), .B2(new_n873), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT121), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n589), .A4(new_n826), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n589), .A3(new_n826), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT122), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n869), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n861), .A2(new_n826), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT59), .B(new_n297), .C1(new_n886), .C2(new_n589), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n868), .B1(new_n885), .B2(new_n887), .ZN(G1345gat));
  NAND3_X1  g687(.A1(new_n867), .A2(new_n305), .A3(new_n511), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n511), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n305), .ZN(G1346gat));
  NAND3_X1  g691(.A1(new_n867), .A2(new_n306), .A3(new_n652), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n886), .A2(new_n652), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(new_n306), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n622), .A2(new_n626), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n789), .B2(new_n791), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n797), .ZN(new_n900));
  AOI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n617), .ZN(new_n901));
  INV_X1    g700(.A(new_n353), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n247), .A3(new_n653), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n904), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n248), .A3(new_n589), .ZN(new_n906));
  OAI21_X1  g705(.A(G176gat), .B1(new_n903), .B2(new_n590), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n900), .A2(new_n217), .A3(new_n511), .ZN(new_n909));
  OAI21_X1  g708(.A(G183gat), .B1(new_n903), .B2(new_n755), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT124), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT123), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n902), .A3(new_n652), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G190gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n919), .B(new_n920), .C1(KEYINPUT126), .C2(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n923), .B(new_n924), .C1(new_n920), .C2(new_n919), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n900), .A2(new_n218), .A3(new_n652), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n643), .A2(new_n898), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n879), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G197gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n653), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n840), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n617), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n931), .A2(new_n934), .ZN(G1352gat));
  NOR3_X1   g734(.A1(new_n932), .A2(G204gat), .A3(new_n590), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n879), .A2(new_n589), .A3(new_n928), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G204gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(G1353gat));
  OAI21_X1  g741(.A(G211gat), .B1(new_n929), .B2(new_n755), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n943), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n944));
  NAND2_X1  g743(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n945));
  OR2_X1    g744(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n933), .A2(new_n314), .A3(new_n511), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(G1354gat));
  OAI21_X1  g748(.A(G218gat), .B1(new_n929), .B2(new_n562), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n315), .A3(new_n652), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1355gat));
endmodule


