

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n696), .A2(n695), .ZN(n704) );
  XNOR2_X1 U553 ( .A(n703), .B(n702), .ZN(n707) );
  INV_X1 U554 ( .A(KEYINPUT99), .ZN(n702) );
  INV_X1 U555 ( .A(n736), .ZN(n697) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n720) );
  XNOR2_X1 U557 ( .A(n721), .B(n720), .ZN(n725) );
  OR2_X1 U558 ( .A1(n751), .A2(n750), .ZN(n767) );
  NAND2_X1 U559 ( .A1(G40), .A2(G160), .ZN(n690) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n640) );
  NOR2_X1 U561 ( .A1(G651), .A2(n653), .ZN(n648) );
  NOR2_X2 U562 ( .A1(n516), .A2(G2104), .ZN(n876) );
  XNOR2_X1 U563 ( .A(n522), .B(n521), .ZN(n881) );
  NOR2_X1 U564 ( .A1(n526), .A2(n525), .ZN(G160) );
  INV_X1 U565 ( .A(G2105), .ZN(n516) );
  NAND2_X1 U566 ( .A1(G125), .A2(n876), .ZN(n517) );
  XNOR2_X1 U567 ( .A(n517), .B(KEYINPUT64), .ZN(n520) );
  AND2_X1 U568 ( .A1(n516), .A2(G2104), .ZN(n880) );
  NAND2_X1 U569 ( .A1(G101), .A2(n880), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n526) );
  XNOR2_X1 U572 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n881), .A2(G137), .ZN(n524) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U576 ( .A1(n877), .A2(G113), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U578 ( .A(KEYINPUT78), .B(KEYINPUT7), .ZN(n541) );
  NAND2_X1 U579 ( .A1(n640), .A2(G89), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n527), .B(KEYINPUT4), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n653) );
  INV_X1 U582 ( .A(G651), .ZN(n531) );
  NOR2_X1 U583 ( .A1(n653), .A2(n531), .ZN(n637) );
  NAND2_X1 U584 ( .A1(G76), .A2(n637), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n530), .B(KEYINPUT5), .ZN(n539) );
  XNOR2_X1 U587 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n537) );
  NOR2_X1 U588 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n532), .Z(n652) );
  NAND2_X1 U590 ( .A1(n652), .A2(G63), .ZN(n533) );
  XNOR2_X1 U591 ( .A(n533), .B(KEYINPUT76), .ZN(n535) );
  NAND2_X1 U592 ( .A1(G51), .A2(n648), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U594 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n541), .B(n540), .ZN(G168) );
  XOR2_X1 U597 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U598 ( .A1(G64), .A2(n652), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G52), .A2(n648), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G90), .A2(n640), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G77), .A2(n637), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U605 ( .A1(n548), .A2(n547), .ZN(G171) );
  INV_X1 U606 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U607 ( .A(G2427), .B(KEYINPUT108), .ZN(n558) );
  XOR2_X1 U608 ( .A(G2443), .B(G2438), .Z(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT107), .B(G2454), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n550), .B(n549), .ZN(n554) );
  XOR2_X1 U611 ( .A(G2430), .B(G2435), .Z(n552) );
  XNOR2_X1 U612 ( .A(G1341), .B(G1348), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U614 ( .A(n554), .B(n553), .Z(n556) );
  XNOR2_X1 U615 ( .A(G2451), .B(G2446), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n558), .B(n557), .ZN(n559) );
  AND2_X1 U618 ( .A1(n559), .A2(G14), .ZN(G401) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U620 ( .A1(G111), .A2(n877), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT82), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G135), .A2(n881), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT81), .B(n561), .Z(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n876), .A2(G123), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT18), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G99), .A2(n880), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n943) );
  XNOR2_X1 U630 ( .A(n943), .B(G2096), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT83), .ZN(n570) );
  OR2_X1 U632 ( .A1(G2100), .A2(n570), .ZN(G156) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G62), .A2(n652), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G50), .A2(n648), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT86), .B(n573), .Z(n577) );
  NAND2_X1 U639 ( .A1(G88), .A2(n640), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G75), .A2(n637), .ZN(n574) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n578) );
  XOR2_X1 U644 ( .A(n578), .B(KEYINPUT10), .Z(n833) );
  NAND2_X1 U645 ( .A1(n833), .A2(G567), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  XNOR2_X1 U647 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G81), .A2(n640), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT68), .ZN(n581) );
  XNOR2_X1 U650 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G68), .A2(n637), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n585), .B(n584), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n652), .A2(G56), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n586), .Z(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT70), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G43), .A2(n648), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n695) );
  INV_X1 U660 ( .A(n695), .ZN(n988) );
  XOR2_X1 U661 ( .A(G860), .B(KEYINPUT71), .Z(n616) );
  NAND2_X1 U662 ( .A1(n988), .A2(n616), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G301), .A2(G868), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT72), .ZN(n603) );
  INV_X1 U665 ( .A(G868), .ZN(n667) );
  NAND2_X1 U666 ( .A1(G79), .A2(n637), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT74), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G66), .A2(n652), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G54), .A2(n648), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G92), .A2(n640), .ZN(n596) );
  XNOR2_X1 U672 ( .A(KEYINPUT73), .B(n596), .ZN(n597) );
  NOR2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U675 ( .A(KEYINPUT15), .B(n601), .Z(n980) );
  NAND2_X1 U676 ( .A1(n667), .A2(n980), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U678 ( .A(KEYINPUT75), .B(n604), .Z(G284) );
  NAND2_X1 U679 ( .A1(G65), .A2(n652), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G53), .A2(n648), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G91), .A2(n640), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G78), .A2(n637), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n716) );
  INV_X1 U686 ( .A(n716), .ZN(G299) );
  NOR2_X1 U687 ( .A1(G286), .A2(n667), .ZN(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT79), .B(n611), .Z(n613) );
  NOR2_X1 U689 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U691 ( .A(KEYINPUT80), .B(n614), .ZN(G297) );
  INV_X1 U692 ( .A(G559), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n980), .A2(n617), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT16), .B(n618), .Z(G148) );
  NOR2_X1 U696 ( .A1(G868), .A2(n695), .ZN(n621) );
  INV_X1 U697 ( .A(n980), .ZN(n705) );
  NAND2_X1 U698 ( .A1(G868), .A2(n705), .ZN(n619) );
  NOR2_X1 U699 ( .A1(G559), .A2(n619), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U701 ( .A1(n705), .A2(G559), .ZN(n664) );
  XOR2_X1 U702 ( .A(n988), .B(n664), .Z(n622) );
  NOR2_X1 U703 ( .A1(n622), .A2(G860), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G67), .A2(n652), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G55), .A2(n648), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G93), .A2(n640), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G80), .A2(n637), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n666) );
  XNOR2_X1 U711 ( .A(n629), .B(n666), .ZN(G145) );
  NAND2_X1 U712 ( .A1(G60), .A2(n652), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G47), .A2(n648), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U715 ( .A(KEYINPUT66), .B(n632), .Z(n636) );
  NAND2_X1 U716 ( .A1(G85), .A2(n640), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G72), .A2(n637), .ZN(n633) );
  AND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G73), .A2(n637), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(KEYINPUT2), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n639), .B(KEYINPUT84), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G86), .A2(n640), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G61), .A2(n652), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G48), .A2(n648), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U729 ( .A(KEYINPUT85), .B(n647), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G49), .A2(n648), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(G288) );
  XOR2_X1 U736 ( .A(G303), .B(G290), .Z(n656) );
  XNOR2_X1 U737 ( .A(n656), .B(G305), .ZN(n660) );
  XNOR2_X1 U738 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U739 ( .A(G288), .B(KEYINPUT87), .ZN(n657) );
  XNOR2_X1 U740 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U741 ( .A(n660), .B(n659), .Z(n662) );
  XOR2_X1 U742 ( .A(G299), .B(n666), .Z(n661) );
  XNOR2_X1 U743 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n663), .B(n988), .ZN(n901) );
  XOR2_X1 U745 ( .A(n901), .B(n664), .Z(n665) );
  NOR2_X1 U746 ( .A1(n667), .A2(n665), .ZN(n669) );
  AND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U748 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U755 ( .A(KEYINPUT67), .B(G132), .ZN(G219) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U758 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G96), .A2(n676), .ZN(n911) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n911), .ZN(n677) );
  XOR2_X1 U761 ( .A(KEYINPUT89), .B(n677), .Z(n681) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U763 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G108), .A2(n679), .ZN(n912) );
  NAND2_X1 U765 ( .A1(G567), .A2(n912), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n681), .A2(n680), .ZN(n858) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n858), .A2(n682), .ZN(n837) );
  NAND2_X1 U769 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G102), .A2(n880), .ZN(n684) );
  NAND2_X1 U771 ( .A1(G138), .A2(n881), .ZN(n683) );
  NAND2_X1 U772 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U773 ( .A1(G126), .A2(n876), .ZN(n686) );
  NAND2_X1 U774 ( .A1(G114), .A2(n877), .ZN(n685) );
  NAND2_X1 U775 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U776 ( .A1(n688), .A2(n687), .ZN(G164) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n783) );
  INV_X1 U778 ( .A(KEYINPUT90), .ZN(n689) );
  XNOR2_X2 U779 ( .A(n690), .B(n689), .ZN(n782) );
  NAND2_X2 U780 ( .A1(n783), .A2(n782), .ZN(n736) );
  NAND2_X1 U781 ( .A1(n697), .A2(G1996), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT26), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G1341), .A2(n736), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n694), .B(KEYINPUT98), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n704), .A2(n705), .ZN(n701) );
  NOR2_X1 U787 ( .A1(G2067), .A2(n736), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n697), .A2(G1348), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n703) );
  OR2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U792 ( .A1(n707), .A2(n706), .ZN(n714) );
  INV_X1 U793 ( .A(G2072), .ZN(n914) );
  NOR2_X1 U794 ( .A1(n736), .A2(n914), .ZN(n709) );
  XNOR2_X1 U795 ( .A(KEYINPUT96), .B(KEYINPUT27), .ZN(n708) );
  XNOR2_X1 U796 ( .A(n709), .B(n708), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n736), .A2(G1956), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U799 ( .A(KEYINPUT97), .B(n712), .ZN(n715) );
  NAND2_X1 U800 ( .A1(n716), .A2(n715), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n719) );
  NOR2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U803 ( .A(n717), .B(KEYINPUT28), .Z(n718) );
  NAND2_X1 U804 ( .A1(n719), .A2(n718), .ZN(n721) );
  OR2_X1 U805 ( .A1(n697), .A2(G1961), .ZN(n723) );
  XNOR2_X1 U806 ( .A(KEYINPUT25), .B(G2078), .ZN(n913) );
  NAND2_X1 U807 ( .A1(n697), .A2(n913), .ZN(n722) );
  NAND2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n731) );
  NAND2_X1 U809 ( .A1(n731), .A2(G171), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n725), .A2(n724), .ZN(n746) );
  NAND2_X1 U811 ( .A1(G8), .A2(n736), .ZN(n777) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n777), .ZN(n748) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n736), .ZN(n747) );
  NOR2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n726) );
  NAND2_X1 U815 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U816 ( .A(KEYINPUT101), .B(n727), .ZN(n729) );
  XOR2_X1 U817 ( .A(KEYINPUT30), .B(KEYINPUT100), .Z(n728) );
  XNOR2_X1 U818 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U819 ( .A1(G168), .A2(n730), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G171), .A2(n731), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n734), .Z(n745) );
  NAND2_X1 U823 ( .A1(n746), .A2(n745), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n735), .A2(G286), .ZN(n742) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n736), .ZN(n737) );
  XNOR2_X1 U826 ( .A(n737), .B(KEYINPUT102), .ZN(n739) );
  NOR2_X1 U827 ( .A1(n777), .A2(G1971), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n740), .A2(G303), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U831 ( .A1(G8), .A2(n743), .ZN(n744) );
  XNOR2_X1 U832 ( .A(n744), .B(KEYINPUT32), .ZN(n768) );
  AND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n751) );
  AND2_X1 U834 ( .A1(G8), .A2(n747), .ZN(n749) );
  OR2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n972) );
  AND2_X1 U837 ( .A1(n767), .A2(n972), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n768), .A2(n752), .ZN(n758) );
  INV_X1 U839 ( .A(n972), .ZN(n754) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n759), .A2(n753), .ZN(n978) );
  OR2_X1 U843 ( .A1(n754), .A2(n978), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n777), .A2(n755), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n766) );
  NAND2_X1 U847 ( .A1(KEYINPUT33), .A2(n759), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n777), .A2(n760), .ZN(n761) );
  XOR2_X1 U849 ( .A(KEYINPUT103), .B(n761), .Z(n764) );
  XOR2_X1 U850 ( .A(G1981), .B(KEYINPUT104), .Z(n762) );
  XNOR2_X1 U851 ( .A(G305), .B(n762), .ZN(n976) );
  INV_X1 U852 ( .A(n976), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  AND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n781) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n771) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n772), .A2(n777), .ZN(n779) );
  XNOR2_X1 U860 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(KEYINPUT94), .ZN(n775) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n775), .B(n774), .ZN(n776) );
  OR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n797) );
  INV_X1 U867 ( .A(n782), .ZN(n784) );
  NOR2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n828) );
  NAND2_X1 U869 ( .A1(G104), .A2(n880), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G140), .A2(n881), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n788) );
  XOR2_X1 U872 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n787) );
  XNOR2_X1 U873 ( .A(n788), .B(n787), .ZN(n793) );
  NAND2_X1 U874 ( .A1(G128), .A2(n876), .ZN(n790) );
  NAND2_X1 U875 ( .A1(G116), .A2(n877), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U877 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U879 ( .A(n794), .B(KEYINPUT36), .ZN(n795) );
  XNOR2_X1 U880 ( .A(n795), .B(KEYINPUT92), .ZN(n898) );
  XNOR2_X1 U881 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U882 ( .A1(n898), .A2(n826), .ZN(n960) );
  NAND2_X1 U883 ( .A1(n828), .A2(n960), .ZN(n824) );
  INV_X1 U884 ( .A(n824), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n813) );
  NAND2_X1 U886 ( .A1(G129), .A2(n876), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G117), .A2(n877), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n880), .A2(G105), .ZN(n800) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n881), .A2(G141), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n889) );
  AND2_X1 U894 ( .A1(n889), .A2(G1996), .ZN(n944) );
  NAND2_X1 U895 ( .A1(G119), .A2(n876), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G107), .A2(n877), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n811) );
  NAND2_X1 U898 ( .A1(G95), .A2(n880), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G131), .A2(n881), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U901 ( .A(KEYINPUT93), .B(n809), .Z(n810) );
  NOR2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n875) );
  INV_X1 U903 ( .A(G1991), .ZN(n838) );
  NOR2_X1 U904 ( .A1(n875), .A2(n838), .ZN(n948) );
  OR2_X1 U905 ( .A1(n944), .A2(n948), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n828), .A2(n812), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n813), .A2(n817), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(KEYINPUT105), .ZN(n816) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U910 ( .A1(n971), .A2(n828), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n831) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n889), .ZN(n938) );
  INV_X1 U913 ( .A(n817), .ZN(n821) );
  AND2_X1 U914 ( .A1(n838), .A2(n875), .ZN(n942) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n818) );
  XNOR2_X1 U916 ( .A(KEYINPUT106), .B(n818), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n942), .A2(n819), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n938), .A2(n822), .ZN(n823) );
  XNOR2_X1 U920 ( .A(KEYINPUT39), .B(n823), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n898), .A2(n826), .ZN(n945) );
  NAND2_X1 U923 ( .A1(n827), .A2(n945), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n833), .ZN(G217) );
  INV_X1 U928 ( .A(n833), .ZN(G223) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT109), .B(n834), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(G661), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G188) );
  XOR2_X1 U934 ( .A(KEYINPUT41), .B(G1986), .Z(n840) );
  XOR2_X1 U935 ( .A(G1996), .B(n838), .Z(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(n841), .B(KEYINPUT112), .Z(n843) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1981), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1956), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U944 ( .A(KEYINPUT111), .B(G2474), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n851) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n853) );
  XOR2_X1 U950 ( .A(G2067), .B(n914), .Z(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U955 ( .A(KEYINPUT110), .B(n858), .Z(G319) );
  NAND2_X1 U956 ( .A1(G124), .A2(n876), .ZN(n859) );
  XOR2_X1 U957 ( .A(KEYINPUT113), .B(n859), .Z(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U959 ( .A1(G112), .A2(n877), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G100), .A2(n880), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G136), .A2(n881), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G103), .A2(n880), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G139), .A2(n881), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U968 ( .A1(n876), .A2(G127), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT115), .B(n869), .Z(n871) );
  NAND2_X1 U970 ( .A1(n877), .A2(G115), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n951) );
  XNOR2_X1 U974 ( .A(n875), .B(n951), .ZN(n897) );
  NAND2_X1 U975 ( .A1(G130), .A2(n876), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G118), .A2(n877), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U978 ( .A1(G106), .A2(n880), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G142), .A2(n881), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  NOR2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n893) );
  XNOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n887), .B(KEYINPUT114), .ZN(n888) );
  XOR2_X1 U985 ( .A(n888), .B(G162), .Z(n891) );
  XOR2_X1 U986 ( .A(G164), .B(n889), .Z(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U988 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U989 ( .A(G160), .B(n943), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U993 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U994 ( .A(n980), .B(G286), .Z(n902) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U996 ( .A(n903), .B(G301), .Z(n904) );
  NOR2_X1 U997 ( .A1(G37), .A2(n904), .ZN(n905) );
  XNOR2_X1 U998 ( .A(KEYINPUT116), .B(n905), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n907), .ZN(n908) );
  AND2_X1 U1002 ( .A1(n908), .A2(G319), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(G225) );
  XNOR2_X1 U1005 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G120), .ZN(G236) );
  INV_X1 U1008 ( .A(G96), .ZN(G221) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(G325) );
  INV_X1 U1011 ( .A(G325), .ZN(G261) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(G303), .ZN(G166) );
  INV_X1 U1014 ( .A(KEYINPUT55), .ZN(n962) );
  XNOR2_X1 U1015 ( .A(G27), .B(n913), .ZN(n925) );
  XOR2_X1 U1016 ( .A(KEYINPUT121), .B(n914), .Z(n915) );
  XNOR2_X1 U1017 ( .A(n915), .B(G33), .ZN(n920) );
  XOR2_X1 U1018 ( .A(G32), .B(G1996), .Z(n916) );
  NAND2_X1 U1019 ( .A1(n916), .A2(G28), .ZN(n918) );
  XNOR2_X1 U1020 ( .A(G26), .B(G2067), .ZN(n917) );
  NOR2_X1 U1021 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G25), .B(G1991), .ZN(n921) );
  XNOR2_X1 U1024 ( .A(KEYINPUT120), .B(n921), .ZN(n922) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n926), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT122), .B(G34), .Z(n928) );
  XNOR2_X1 U1029 ( .A(G2084), .B(KEYINPUT54), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(n928), .B(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G35), .B(G2090), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1034 ( .A(n962), .B(n933), .Z(n935) );
  INV_X1 U1035 ( .A(G29), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n936), .A2(G11), .ZN(n967) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1040 ( .A(KEYINPUT118), .B(n939), .Z(n940) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n958) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G2084), .B(G160), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n956) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n953) );
  XOR2_X1 U1049 ( .A(G2072), .B(n951), .Z(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1051 ( .A(KEYINPUT50), .B(n954), .Z(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT52), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(G29), .A2(n964), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT119), .B(n965), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n994) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XOR2_X1 U1061 ( .A(G299), .B(G1956), .Z(n969) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n987) );
  XOR2_X1 U1066 ( .A(G1966), .B(KEYINPUT123), .Z(n974) );
  XNOR2_X1 U1067 ( .A(G168), .B(n974), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(KEYINPUT57), .ZN(n985) );
  XOR2_X1 U1070 ( .A(G301), .B(G1961), .Z(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G1348), .B(n980), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G1341), .B(n988), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G1966), .B(G21), .Z(n1004) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n995), .B(G4), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G20), .B(G1956), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(n1002), .B(KEYINPUT60), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(n1005), .B(KEYINPUT125), .ZN(n1013) );
  XOR2_X1 U1093 ( .A(G1986), .B(KEYINPUT126), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(G24), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1971), .B(G22), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G23), .B(G1976), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1011), .Z(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G5), .B(G1961), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1016), .Z(n1017) );
  NOR2_X1 U1104 ( .A1(G16), .A2(n1017), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1018), .Z(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

