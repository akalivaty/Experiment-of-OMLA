

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XOR2_X2 U322 ( .A(n366), .B(n365), .Z(n575) );
  NOR2_X1 U323 ( .A1(n541), .A2(n518), .ZN(n431) );
  XNOR2_X1 U324 ( .A(n418), .B(n417), .ZN(n541) );
  INV_X1 U325 ( .A(n424), .ZN(n400) );
  XNOR2_X1 U326 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U327 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U328 ( .A(n480), .B(n409), .Z(n558) );
  NOR2_X1 U329 ( .A1(n521), .A2(n456), .ZN(n563) );
  XNOR2_X1 U330 ( .A(n458), .B(G190GAT), .ZN(n459) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G176GAT), .B(G183GAT), .Z(n291) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U335 ( .A(KEYINPUT92), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U338 ( .A(n295), .B(n294), .Z(n430) );
  XNOR2_X1 U339 ( .A(G99GAT), .B(G71GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n296), .B(G120GAT), .ZN(n394) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n297), .B(KEYINPUT88), .ZN(n441) );
  XNOR2_X1 U343 ( .A(n394), .B(n441), .ZN(n307) );
  XOR2_X1 U344 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U345 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U347 ( .A(KEYINPUT91), .B(KEYINPUT65), .Z(n301) );
  XOR2_X1 U348 ( .A(G43GAT), .B(G134GAT), .Z(n384) );
  XOR2_X1 U349 ( .A(G15GAT), .B(G127GAT), .Z(n353) );
  XNOR2_X1 U350 ( .A(n384), .B(n353), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(n303), .B(n302), .Z(n305) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n430), .B(n308), .Z(n531) );
  INV_X1 U357 ( .A(n531), .ZN(n521) );
  XOR2_X1 U358 ( .A(G78GAT), .B(G148GAT), .Z(n310) );
  XNOR2_X1 U359 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n393) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G162GAT), .Z(n380) );
  XOR2_X1 U362 ( .A(n393), .B(n380), .Z(n312) );
  NAND2_X1 U363 ( .A1(G228GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n324) );
  XOR2_X1 U365 ( .A(G204GAT), .B(KEYINPUT98), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT99), .B(KEYINPUT95), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U368 ( .A(n315), .B(KEYINPUT100), .Z(n317) );
  XOR2_X1 U369 ( .A(G22GAT), .B(G155GAT), .Z(n349) );
  XNOR2_X1 U370 ( .A(n349), .B(KEYINPUT22), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n318), .B(KEYINPUT24), .Z(n322) );
  XOR2_X1 U373 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n320) );
  XNOR2_X1 U374 ( .A(G141GAT), .B(KEYINPUT97), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n440) );
  XNOR2_X1 U376 ( .A(n440), .B(KEYINPUT23), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT96), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U380 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U382 ( .A(G197GAT), .B(n327), .Z(n422) );
  XOR2_X1 U383 ( .A(n328), .B(n422), .Z(n470) );
  XOR2_X1 U384 ( .A(G113GAT), .B(G36GAT), .Z(n330) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G50GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U387 ( .A(n331), .B(G15GAT), .Z(n333) );
  XOR2_X1 U388 ( .A(G1GAT), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(n354), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n334), .B(KEYINPUT8), .ZN(n370) );
  XOR2_X1 U393 ( .A(n370), .B(KEYINPUT68), .Z(n336) );
  NAND2_X1 U394 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(n338), .B(n337), .Z(n346) );
  XOR2_X1 U397 ( .A(KEYINPUT71), .B(G197GAT), .Z(n340) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(G22GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n342) );
  XNOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(n346), .B(n345), .Z(n544) );
  INV_X1 U405 ( .A(n544), .ZN(n568) );
  XOR2_X1 U406 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n348) );
  XNOR2_X1 U407 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n366) );
  XOR2_X1 U409 ( .A(n349), .B(KEYINPUT85), .Z(n351) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n364) );
  XOR2_X1 U413 ( .A(G57GAT), .B(KEYINPUT13), .Z(n397) );
  XOR2_X1 U414 ( .A(n397), .B(G78GAT), .Z(n356) );
  XNOR2_X1 U415 ( .A(n354), .B(G211GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U417 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT84), .B(KEYINPUT14), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U420 ( .A(n360), .B(n359), .Z(n362) );
  XNOR2_X1 U421 ( .A(G183GAT), .B(G71GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  INV_X1 U424 ( .A(n575), .ZN(n551) );
  XOR2_X1 U425 ( .A(KEYINPUT66), .B(KEYINPUT77), .Z(n372) );
  XOR2_X1 U426 ( .A(KEYINPUT10), .B(G106GAT), .Z(n368) );
  XNOR2_X1 U427 ( .A(G190GAT), .B(G99GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n379) );
  XOR2_X1 U431 ( .A(KEYINPUT9), .B(KEYINPUT67), .Z(n374) );
  XNOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT11), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U434 ( .A(n375), .B(KEYINPUT78), .Z(n377) );
  XOR2_X1 U435 ( .A(G85GAT), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U436 ( .A(G218GAT), .B(n398), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(n379), .B(n378), .Z(n386) );
  XOR2_X1 U439 ( .A(G36GAT), .B(KEYINPUT80), .Z(n423) );
  XOR2_X1 U440 ( .A(n380), .B(n423), .Z(n382) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n457) );
  XOR2_X1 U445 ( .A(n457), .B(KEYINPUT36), .Z(n579) );
  NOR2_X1 U446 ( .A1(n551), .A2(n579), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n387), .B(KEYINPUT45), .ZN(n406) );
  XOR2_X1 U448 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n389) );
  XNOR2_X1 U449 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n388) );
  XOR2_X1 U450 ( .A(n389), .B(n388), .Z(n405) );
  XOR2_X1 U451 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n391) );
  NAND2_X1 U452 ( .A1(G230GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U454 ( .A(n392), .B(KEYINPUT72), .Z(n396) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n401) );
  XNOR2_X1 U458 ( .A(G204GAT), .B(G64GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n399), .B(KEYINPUT76), .ZN(n424) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n572) );
  INV_X1 U461 ( .A(n572), .ZN(n480) );
  NAND2_X1 U462 ( .A1(n406), .A2(n480), .ZN(n407) );
  NOR2_X1 U463 ( .A1(n568), .A2(n407), .ZN(n408) );
  XOR2_X1 U464 ( .A(KEYINPUT120), .B(n408), .Z(n416) );
  XOR2_X1 U465 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n409) );
  NAND2_X1 U466 ( .A1(n568), .A2(n558), .ZN(n410) );
  XOR2_X1 U467 ( .A(KEYINPUT46), .B(n410), .Z(n411) );
  NOR2_X1 U468 ( .A1(n575), .A2(n411), .ZN(n412) );
  INV_X1 U469 ( .A(n457), .ZN(n554) );
  NAND2_X1 U470 ( .A1(n412), .A2(n554), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n413), .B(KEYINPUT119), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n414), .B(KEYINPUT47), .ZN(n415) );
  NAND2_X1 U473 ( .A1(n416), .A2(n415), .ZN(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT121), .B(KEYINPUT48), .ZN(n417) );
  XOR2_X1 U475 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n420) );
  XNOR2_X1 U476 ( .A(G8GAT), .B(G92GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U479 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U480 ( .A1(G226GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n518) );
  XNOR2_X1 U484 ( .A(n431), .B(KEYINPUT54), .ZN(n454) );
  XOR2_X1 U485 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n433) );
  XNOR2_X1 U486 ( .A(KEYINPUT4), .B(KEYINPUT103), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n445) );
  XOR2_X1 U488 ( .A(KEYINPUT101), .B(G155GAT), .Z(n435) );
  XNOR2_X1 U489 ( .A(G127GAT), .B(G148GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U491 ( .A(G57GAT), .B(KEYINPUT5), .Z(n437) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n453) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n451) );
  XOR2_X1 U499 ( .A(G85GAT), .B(G162GAT), .Z(n447) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(G134GAT), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U502 ( .A(G29GAT), .B(KEYINPUT79), .Z(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n516) );
  NAND2_X1 U506 ( .A1(n454), .A2(n516), .ZN(n566) );
  NOR2_X1 U507 ( .A1(n470), .A2(n566), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NAND2_X1 U509 ( .A1(n563), .A2(n457), .ZN(n460) );
  XOR2_X1 U510 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n458) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n518), .ZN(n469) );
  NAND2_X1 U512 ( .A1(n470), .A2(n521), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(KEYINPUT26), .ZN(n567) );
  NOR2_X1 U514 ( .A1(n469), .A2(n567), .ZN(n462) );
  XNOR2_X1 U515 ( .A(KEYINPUT107), .B(n462), .ZN(n466) );
  NOR2_X1 U516 ( .A1(n521), .A2(n518), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n470), .A2(n463), .ZN(n464) );
  XNOR2_X1 U518 ( .A(KEYINPUT25), .B(n464), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n516), .A2(n467), .ZN(n468) );
  XOR2_X1 U521 ( .A(KEYINPUT108), .B(n468), .Z(n474) );
  NOR2_X1 U522 ( .A1(n469), .A2(n516), .ZN(n543) );
  XOR2_X1 U523 ( .A(KEYINPUT28), .B(n470), .Z(n525) );
  NAND2_X1 U524 ( .A1(n543), .A2(n525), .ZN(n529) );
  XNOR2_X1 U525 ( .A(KEYINPUT94), .B(n531), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n529), .A2(n471), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT106), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n474), .A2(n473), .ZN(n490) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(KEYINPUT87), .Z(n476) );
  NAND2_X1 U530 ( .A1(n575), .A2(n554), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U532 ( .A(n477), .B(KEYINPUT86), .ZN(n478) );
  NOR2_X1 U533 ( .A1(n490), .A2(n478), .ZN(n479) );
  XNOR2_X1 U534 ( .A(KEYINPUT109), .B(n479), .ZN(n504) );
  NAND2_X1 U535 ( .A1(n568), .A2(n480), .ZN(n494) );
  NOR2_X1 U536 ( .A1(n504), .A2(n494), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT110), .B(n481), .Z(n488) );
  NOR2_X1 U538 ( .A1(n488), .A2(n516), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT34), .B(n482), .Z(n483) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n488), .A2(n518), .ZN(n484) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n484), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n488), .A2(n521), .ZN(n486) );
  XNOR2_X1 U544 ( .A(KEYINPUT111), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  NOR2_X1 U547 ( .A1(n488), .A2(n525), .ZN(n489) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT112), .B(KEYINPUT37), .Z(n493) );
  NOR2_X1 U550 ( .A1(n490), .A2(n579), .ZN(n491) );
  NAND2_X1 U551 ( .A1(n491), .A2(n551), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n515) );
  NOR2_X1 U553 ( .A1(n515), .A2(n494), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n495), .Z(n502) );
  NOR2_X1 U555 ( .A1(n502), .A2(n516), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n502), .A2(n518), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT113), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1329GAT) );
  NOR2_X1 U561 ( .A1(n502), .A2(n521), .ZN(n500) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n502), .A2(n525), .ZN(n503) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  NAND2_X1 U566 ( .A1(n544), .A2(n558), .ZN(n514) );
  OR2_X1 U567 ( .A1(n504), .A2(n514), .ZN(n511) );
  NOR2_X1 U568 ( .A1(n516), .A2(n511), .ZN(n506) );
  XNOR2_X1 U569 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n507), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n518), .A2(n511), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(KEYINPUT115), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U575 ( .A1(n521), .A2(n511), .ZN(n510) );
  XOR2_X1 U576 ( .A(G71GAT), .B(n510), .Z(G1334GAT) );
  NOR2_X1 U577 ( .A1(n525), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  OR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n516), .A2(n524), .ZN(n517) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n524), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT116), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n524), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT117), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT118), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n541), .A2(n529), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n544), .A2(n537), .ZN(n532) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  INV_X1 U597 ( .A(n558), .ZN(n546) );
  NOR2_X1 U598 ( .A1(n546), .A2(n537), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n551), .A2(n537), .ZN(n535) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(n535), .Z(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n554), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT122), .B(KEYINPUT51), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n567), .A2(n541), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n544), .A2(n553), .ZN(n545) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n553), .A2(n546), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT123), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT124), .B(n555), .Z(n556) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n563), .A2(n568), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n560) );
  NAND2_X1 U625 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n575), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT126), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(n565), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n577), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n577), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U642 ( .A(n577), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

