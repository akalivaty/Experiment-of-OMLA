

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n318) );
  XNOR2_X1 U325 ( .A(n473), .B(n472), .ZN(n478) );
  XNOR2_X1 U326 ( .A(n487), .B(n486), .ZN(n525) );
  XOR2_X1 U327 ( .A(n347), .B(KEYINPUT7), .Z(n292) );
  XNOR2_X1 U328 ( .A(n471), .B(KEYINPUT25), .ZN(n472) );
  INV_X1 U329 ( .A(KEYINPUT18), .ZN(n319) );
  XNOR2_X1 U330 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U331 ( .A(n322), .B(n321), .ZN(n445) );
  NOR2_X1 U332 ( .A1(n480), .A2(n495), .ZN(n481) );
  XNOR2_X1 U333 ( .A(n305), .B(n304), .ZN(n306) );
  NOR2_X1 U334 ( .A1(n422), .A2(n495), .ZN(n577) );
  XNOR2_X1 U335 ( .A(n307), .B(n306), .ZN(n312) );
  XNOR2_X1 U336 ( .A(n398), .B(KEYINPUT48), .ZN(n555) );
  XOR2_X1 U337 ( .A(n435), .B(n333), .Z(n468) );
  INV_X1 U338 ( .A(KEYINPUT58), .ZN(n461) );
  XNOR2_X1 U339 ( .A(n461), .B(G190GAT), .ZN(n462) );
  XNOR2_X1 U340 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(G85GAT), .B(G99GAT), .Z(n338) );
  XOR2_X1 U342 ( .A(G64GAT), .B(G204GAT), .Z(n331) );
  XOR2_X1 U343 ( .A(G120GAT), .B(G71GAT), .Z(n451) );
  XOR2_X1 U344 ( .A(n331), .B(n451), .Z(n294) );
  NAND2_X1 U345 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n338), .B(n295), .ZN(n307) );
  XOR2_X1 U348 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n297) );
  XNOR2_X1 U349 ( .A(G92GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT76), .B(KEYINPUT79), .Z(n299) );
  XNOR2_X1 U352 ( .A(KEYINPUT80), .B(KEYINPUT74), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(n301), .B(n300), .Z(n305) );
  XOR2_X1 U355 ( .A(KEYINPUT32), .B(KEYINPUT78), .Z(n303) );
  XNOR2_X1 U356 ( .A(KEYINPUT31), .B(KEYINPUT75), .ZN(n302) );
  XOR2_X1 U357 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U358 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n308), .B(KEYINPUT72), .ZN(n376) );
  XOR2_X1 U360 ( .A(KEYINPUT77), .B(G78GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(G148GAT), .B(G106GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n426) );
  XNOR2_X1 U363 ( .A(n376), .B(n426), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n583) );
  XNOR2_X1 U365 ( .A(n583), .B(KEYINPUT41), .ZN(n544) );
  XOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT92), .Z(n314) );
  XNOR2_X1 U367 ( .A(KEYINPUT93), .B(KEYINPUT21), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n315), .B(KEYINPUT94), .Z(n317) );
  XNOR2_X1 U370 ( .A(G218GAT), .B(G211GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n435) );
  XNOR2_X1 U372 ( .A(n318), .B(G176GAT), .ZN(n322) );
  XNOR2_X1 U373 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n320) );
  XOR2_X1 U374 ( .A(G190GAT), .B(G92GAT), .Z(n349) );
  XNOR2_X1 U375 ( .A(n445), .B(n349), .ZN(n326) );
  INV_X1 U376 ( .A(n326), .ZN(n324) );
  AND2_X1 U377 ( .A1(G226GAT), .A2(G233GAT), .ZN(n325) );
  INV_X1 U378 ( .A(n325), .ZN(n323) );
  NAND2_X1 U379 ( .A1(n324), .A2(n323), .ZN(n328) );
  NAND2_X1 U380 ( .A1(n326), .A2(n325), .ZN(n327) );
  NAND2_X1 U381 ( .A1(n328), .A2(n327), .ZN(n330) );
  XOR2_X1 U382 ( .A(G36GAT), .B(G8GAT), .Z(n329) );
  XOR2_X1 U383 ( .A(G169GAT), .B(n329), .Z(n357) );
  XNOR2_X1 U384 ( .A(n330), .B(n357), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  INV_X1 U386 ( .A(n468), .ZN(n528) );
  XOR2_X1 U387 ( .A(n528), .B(KEYINPUT120), .Z(n399) );
  XOR2_X1 U388 ( .A(KEYINPUT82), .B(KEYINPUT9), .Z(n335) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(G36GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n353) );
  XOR2_X1 U391 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n337) );
  XNOR2_X1 U392 ( .A(G218GAT), .B(KEYINPUT83), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n339) );
  XOR2_X1 U394 ( .A(n339), .B(n338), .Z(n341) );
  XNOR2_X1 U395 ( .A(G162GAT), .B(G134GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U397 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n343) );
  NAND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n351) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(KEYINPUT70), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n346), .B(KEYINPUT8), .ZN(n347) );
  XNOR2_X1 U403 ( .A(G29GAT), .B(G43GAT), .ZN(n348) );
  XOR2_X1 U404 ( .A(n292), .B(n348), .Z(n367) );
  XNOR2_X1 U405 ( .A(n367), .B(n349), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X2 U407 ( .A(n353), .B(n352), .Z(n551) );
  INV_X1 U408 ( .A(n551), .ZN(n568) );
  INV_X1 U409 ( .A(n544), .ZN(n561) );
  XOR2_X1 U410 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n355) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U412 ( .A(G113GAT), .B(G15GAT), .Z(n448) );
  XNOR2_X1 U413 ( .A(n431), .B(n448), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n356), .B(KEYINPUT65), .Z(n362) );
  XOR2_X1 U416 ( .A(n357), .B(KEYINPUT66), .Z(n359) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(n360), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n364) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(KEYINPUT29), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n580) );
  NAND2_X1 U426 ( .A1(n561), .A2(n580), .ZN(n369) );
  XNOR2_X1 U427 ( .A(KEYINPUT46), .B(n369), .ZN(n389) );
  XOR2_X1 U428 ( .A(KEYINPUT84), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U429 ( .A(G1GAT), .B(G8GAT), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT86), .B(KEYINPUT12), .Z(n373) );
  XNOR2_X1 U432 ( .A(KEYINPUT15), .B(KEYINPUT85), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n388) );
  XOR2_X1 U435 ( .A(n376), .B(KEYINPUT14), .Z(n378) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U438 ( .A(G15GAT), .B(G71GAT), .Z(n380) );
  XNOR2_X1 U439 ( .A(G127GAT), .B(G183GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U442 ( .A(G211GAT), .B(G22GAT), .Z(n384) );
  XNOR2_X1 U443 ( .A(G155GAT), .B(G78GAT), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U446 ( .A(n388), .B(n387), .Z(n587) );
  INV_X1 U447 ( .A(n587), .ZN(n573) );
  NAND2_X1 U448 ( .A1(n389), .A2(n573), .ZN(n390) );
  NOR2_X1 U449 ( .A1(n568), .A2(n390), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT47), .ZN(n397) );
  XOR2_X1 U451 ( .A(KEYINPUT36), .B(n551), .Z(n589) );
  AND2_X1 U452 ( .A1(n589), .A2(n587), .ZN(n393) );
  INV_X1 U453 ( .A(KEYINPUT45), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n394) );
  NOR2_X1 U455 ( .A1(n583), .A2(n394), .ZN(n395) );
  XNOR2_X1 U456 ( .A(KEYINPUT71), .B(n580), .ZN(n541) );
  NAND2_X1 U457 ( .A1(n395), .A2(n541), .ZN(n396) );
  NAND2_X1 U458 ( .A1(n397), .A2(n396), .ZN(n398) );
  NAND2_X1 U459 ( .A1(n399), .A2(n555), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT54), .ZN(n401) );
  XOR2_X1 U461 ( .A(KEYINPUT121), .B(n401), .Z(n422) );
  XOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT95), .Z(n403) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G57GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n421) );
  XOR2_X1 U465 ( .A(G113GAT), .B(G120GAT), .Z(n405) );
  XNOR2_X1 U466 ( .A(G148GAT), .B(G141GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U468 ( .A(G29GAT), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n417) );
  XOR2_X1 U470 ( .A(G155GAT), .B(KEYINPUT2), .Z(n409) );
  XNOR2_X1 U471 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n427) );
  XOR2_X1 U473 ( .A(G127GAT), .B(KEYINPUT0), .Z(n411) );
  XNOR2_X1 U474 ( .A(G134GAT), .B(KEYINPUT87), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n450) );
  XNOR2_X1 U476 ( .A(n427), .B(n450), .ZN(n415) );
  XOR2_X1 U477 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n413) );
  XNOR2_X1 U478 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n419) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n495) );
  XOR2_X1 U485 ( .A(G204GAT), .B(KEYINPUT22), .Z(n424) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U488 ( .A(n425), .B(KEYINPUT24), .Z(n429) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U491 ( .A(n430), .B(KEYINPUT23), .Z(n433) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n474) );
  NAND2_X1 U495 ( .A1(n577), .A2(n474), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n436) );
  XNOR2_X1 U497 ( .A(KEYINPUT55), .B(n436), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n454) );
  XOR2_X1 U499 ( .A(KEYINPUT20), .B(G169GAT), .Z(n440) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(n441), .B(KEYINPUT89), .Z(n447) );
  XOR2_X1 U503 ( .A(KEYINPUT88), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G190GAT), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n453) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U510 ( .A(n453), .B(n452), .Z(n469) );
  NAND2_X1 U511 ( .A1(n454), .A2(n469), .ZN(n572) );
  NOR2_X1 U512 ( .A1(n544), .A2(n572), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(G176GAT), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  NOR2_X1 U516 ( .A1(n541), .A2(n572), .ZN(n460) );
  INV_X1 U517 ( .A(G169GAT), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n458), .B(KEYINPUT124), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(G1348GAT) );
  NOR2_X1 U520 ( .A1(n551), .A2(n572), .ZN(n463) );
  INV_X1 U521 ( .A(G43GAT), .ZN(n492) );
  INV_X1 U522 ( .A(n469), .ZN(n539) );
  XOR2_X1 U523 ( .A(KEYINPUT107), .B(KEYINPUT38), .Z(n489) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n464) );
  XOR2_X1 U525 ( .A(n468), .B(n464), .Z(n477) );
  XOR2_X1 U526 ( .A(KEYINPUT28), .B(n474), .Z(n506) );
  NOR2_X1 U527 ( .A1(n477), .A2(n506), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n465), .A2(n495), .ZN(n538) );
  XOR2_X1 U529 ( .A(KEYINPUT91), .B(n469), .Z(n466) );
  NOR2_X1 U530 ( .A1(n538), .A2(n466), .ZN(n467) );
  XOR2_X1 U531 ( .A(KEYINPUT98), .B(n467), .Z(n483) );
  NAND2_X1 U532 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U533 ( .A1(n470), .A2(n474), .ZN(n473) );
  INV_X1 U534 ( .A(KEYINPUT99), .ZN(n471) );
  INV_X1 U535 ( .A(n474), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n539), .A2(n475), .ZN(n476) );
  XNOR2_X1 U537 ( .A(KEYINPUT26), .B(n476), .ZN(n579) );
  NOR2_X1 U538 ( .A1(n579), .A2(n477), .ZN(n556) );
  NOR2_X1 U539 ( .A1(n478), .A2(n556), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT100), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT101), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n498) );
  NAND2_X1 U543 ( .A1(n498), .A2(n573), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT105), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n485), .A2(n589), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n486) );
  NOR2_X1 U547 ( .A1(n583), .A2(n541), .ZN(n499) );
  NAND2_X1 U548 ( .A1(n525), .A2(n499), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n513) );
  NOR2_X1 U550 ( .A1(n539), .A2(n513), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1330GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n494) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n501) );
  INV_X1 U556 ( .A(n495), .ZN(n557) );
  NAND2_X1 U557 ( .A1(n551), .A2(n587), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT16), .B(n496), .Z(n497) );
  AND2_X1 U559 ( .A1(n498), .A2(n497), .ZN(n516) );
  NAND2_X1 U560 ( .A1(n499), .A2(n516), .ZN(n507) );
  NOR2_X1 U561 ( .A1(n557), .A2(n507), .ZN(n500) );
  XOR2_X1 U562 ( .A(n501), .B(n500), .Z(G1324GAT) );
  NOR2_X1 U563 ( .A1(n528), .A2(n507), .ZN(n502) );
  XOR2_X1 U564 ( .A(G8GAT), .B(n502), .Z(G1325GAT) );
  NOR2_X1 U565 ( .A1(n539), .A2(n507), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G15GAT), .B(n505), .ZN(G1326GAT) );
  INV_X1 U569 ( .A(n506), .ZN(n535) );
  NOR2_X1 U570 ( .A1(n535), .A2(n507), .ZN(n508) );
  XOR2_X1 U571 ( .A(G22GAT), .B(n508), .Z(G1327GAT) );
  NOR2_X1 U572 ( .A1(n557), .A2(n513), .ZN(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT39), .B(KEYINPUT108), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G29GAT), .ZN(G1328GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n528), .ZN(n512) );
  XOR2_X1 U577 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n535), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  NOR2_X1 U581 ( .A1(n544), .A2(n580), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n526), .A2(n516), .ZN(n522) );
  NOR2_X1 U583 ( .A1(n557), .A2(n522), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U586 ( .A(G57GAT), .B(n519), .Z(G1332GAT) );
  NOR2_X1 U587 ( .A1(n528), .A2(n522), .ZN(n520) );
  XOR2_X1 U588 ( .A(G64GAT), .B(n520), .Z(G1333GAT) );
  NOR2_X1 U589 ( .A1(n539), .A2(n522), .ZN(n521) );
  XOR2_X1 U590 ( .A(G71GAT), .B(n521), .Z(G1334GAT) );
  NOR2_X1 U591 ( .A1(n535), .A2(n522), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n534) );
  NOR2_X1 U595 ( .A1(n557), .A2(n534), .ZN(n527) );
  XOR2_X1 U596 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U597 ( .A1(n528), .A2(n534), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(G1337GAT) );
  INV_X1 U600 ( .A(KEYINPUT112), .ZN(n532) );
  NOR2_X1 U601 ( .A1(n539), .A2(n534), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U603 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U605 ( .A(KEYINPUT44), .B(n536), .Z(n537) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U608 ( .A1(n555), .A2(n540), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n541), .A2(n550), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n550), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NOR2_X1 U615 ( .A1(n573), .A2(n550), .ZN(n548) );
  XNOR2_X1 U616 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U618 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U620 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(G134GAT), .B(n554), .Z(G1343GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT116), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n569), .A2(n580), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n563) );
  NAND2_X1 U629 ( .A1(n561), .A2(n569), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT53), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n587), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT118), .ZN(n567) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n567), .ZN(G1346GAT) );
  XOR2_X1 U636 ( .A(G162GAT), .B(KEYINPUT119), .Z(n571) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1347GAT) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n582) );
  INV_X1 U644 ( .A(n577), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n580), .A2(n590), .ZN(n581) );
  XOR2_X1 U647 ( .A(n582), .B(n581), .Z(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n590), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n590), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U654 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n592) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

