

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761;

  XNOR2_X1 U370 ( .A(n388), .B(G119), .ZN(n390) );
  INV_X1 U371 ( .A(G146), .ZN(n387) );
  OR2_X2 U372 ( .A1(n366), .A2(KEYINPUT53), .ZN(n355) );
  XNOR2_X1 U373 ( .A(n499), .B(n498), .ZN(n504) );
  XNOR2_X2 U374 ( .A(n444), .B(n443), .ZN(n577) );
  XOR2_X2 U375 ( .A(KEYINPUT42), .B(n555), .Z(n760) );
  AND2_X2 U376 ( .A1(n504), .A2(n559), .ZN(n511) );
  XNOR2_X2 U377 ( .A(n558), .B(n557), .ZN(n732) );
  XNOR2_X2 U378 ( .A(n503), .B(KEYINPUT32), .ZN(n636) );
  XNOR2_X2 U379 ( .A(n745), .B(n437), .ZN(n620) );
  XNOR2_X2 U380 ( .A(n432), .B(n385), .ZN(n480) );
  XNOR2_X2 U381 ( .A(n384), .B(G128), .ZN(n432) );
  XNOR2_X2 U382 ( .A(n428), .B(n427), .ZN(n745) );
  XOR2_X2 U383 ( .A(n553), .B(n552), .Z(n684) );
  NOR2_X2 U384 ( .A1(n655), .A2(n656), .ZN(n553) );
  XNOR2_X1 U385 ( .A(n359), .B(n414), .ZN(n374) );
  INV_X2 U386 ( .A(G953), .ZN(n756) );
  NAND2_X1 U387 ( .A1(n357), .A2(n378), .ZN(n513) );
  NOR2_X1 U388 ( .A1(n598), .A2(n601), .ZN(n566) );
  NAND2_X1 U389 ( .A1(n516), .A2(n515), .ZN(n514) );
  XNOR2_X1 U390 ( .A(n375), .B(n374), .ZN(n373) );
  AND2_X1 U391 ( .A1(n365), .A2(n355), .ZN(n364) );
  NAND2_X1 U392 ( .A1(n361), .A2(n368), .ZN(n367) );
  NAND2_X1 U393 ( .A1(n609), .A2(n608), .ZN(n628) );
  AND2_X1 U394 ( .A1(n521), .A2(n549), .ZN(n539) );
  AND2_X1 U395 ( .A1(n500), .A2(n663), .ZN(n521) );
  XNOR2_X1 U396 ( .A(n373), .B(n750), .ZN(n699) );
  INV_X2 U397 ( .A(KEYINPUT3), .ZN(n388) );
  INV_X1 U398 ( .A(G143), .ZN(n384) );
  INV_X1 U399 ( .A(n640), .ZN(n610) );
  AND2_X1 U400 ( .A1(n628), .A2(n349), .ZN(n622) );
  AND2_X1 U401 ( .A1(n627), .A2(G210), .ZN(n349) );
  INV_X1 U402 ( .A(n618), .ZN(n350) );
  AND2_X2 U403 ( .A1(n628), .A2(n627), .ZN(n707) );
  OR2_X2 U404 ( .A1(n640), .A2(KEYINPUT75), .ZN(n641) );
  INV_X1 U405 ( .A(n610), .ZN(n351) );
  INV_X1 U406 ( .A(n351), .ZN(n352) );
  XNOR2_X2 U407 ( .A(n353), .B(n354), .ZN(n565) );
  NOR2_X1 U408 ( .A1(n620), .A2(n531), .ZN(n353) );
  NOR2_X1 U409 ( .A1(n441), .A2(n617), .ZN(n354) );
  XNOR2_X2 U410 ( .A(n530), .B(n529), .ZN(n640) );
  AND2_X2 U411 ( .A1(n692), .A2(n525), .ZN(n381) );
  XNOR2_X2 U412 ( .A(n513), .B(KEYINPUT106), .ZN(n692) );
  OR2_X1 U413 ( .A1(n689), .A2(n371), .ZN(n370) );
  INV_X1 U414 ( .A(KEYINPUT110), .ZN(n538) );
  XNOR2_X1 U415 ( .A(n377), .B(n376), .ZN(n597) );
  INV_X1 U416 ( .A(KEYINPUT39), .ZN(n376) );
  NAND2_X1 U417 ( .A1(n667), .A2(n360), .ZN(n668) );
  INV_X1 U418 ( .A(n521), .ZN(n360) );
  XNOR2_X1 U419 ( .A(KEYINPUT48), .B(KEYINPUT79), .ZN(n595) );
  XNOR2_X1 U420 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U421 ( .A(n383), .B(n433), .ZN(n386) );
  OR2_X2 U422 ( .A1(n710), .A2(G902), .ZN(n404) );
  AND2_X1 U423 ( .A1(n369), .A2(n756), .ZN(n368) );
  NAND2_X1 U424 ( .A1(n689), .A2(n371), .ZN(n369) );
  NOR2_X1 U425 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U426 ( .A1(n732), .A2(n652), .ZN(n563) );
  OR2_X1 U427 ( .A1(n683), .A2(n493), .ZN(n458) );
  AND2_X1 U428 ( .A1(n543), .A2(n542), .ZN(n571) );
  AND2_X1 U429 ( .A1(n366), .A2(KEYINPUT53), .ZN(n356) );
  XOR2_X1 U430 ( .A(n512), .B(KEYINPUT80), .Z(n357) );
  XNOR2_X1 U431 ( .A(n549), .B(KEYINPUT1), .ZN(n501) );
  XOR2_X1 U432 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n358) );
  XOR2_X1 U433 ( .A(n411), .B(n358), .Z(n359) );
  INV_X1 U434 ( .A(KEYINPUT53), .ZN(n372) );
  XNOR2_X2 U435 ( .A(n456), .B(n455), .ZN(n493) );
  OR2_X1 U436 ( .A1(n690), .A2(n370), .ZN(n361) );
  NAND2_X1 U437 ( .A1(n364), .A2(n362), .ZN(G75) );
  NAND2_X1 U438 ( .A1(n363), .A2(n356), .ZN(n362) );
  INV_X1 U439 ( .A(n367), .ZN(n363) );
  NAND2_X1 U440 ( .A1(n367), .A2(n372), .ZN(n365) );
  NAND2_X1 U441 ( .A1(n690), .A2(n371), .ZN(n366) );
  INV_X1 U442 ( .A(KEYINPUT123), .ZN(n371) );
  NAND2_X1 U443 ( .A1(n699), .A2(n486), .ZN(n420) );
  NAND2_X1 U444 ( .A1(n481), .A2(G221), .ZN(n375) );
  NOR2_X1 U445 ( .A1(n597), .A2(n558), .ZN(n544) );
  NAND2_X1 U446 ( .A1(n571), .A2(n653), .ZN(n377) );
  BUF_X1 U447 ( .A(n500), .Z(n662) );
  XNOR2_X2 U448 ( .A(KEYINPUT105), .B(n518), .ZN(n657) );
  XNOR2_X1 U449 ( .A(n420), .B(n419), .ZN(n500) );
  XNOR2_X1 U450 ( .A(n539), .B(n538), .ZN(n540) );
  NOR2_X1 U451 ( .A1(n647), .A2(n352), .ZN(n648) );
  AND2_X1 U452 ( .A1(n662), .A2(n667), .ZN(n378) );
  NOR2_X1 U453 ( .A1(n655), .A2(n495), .ZN(n379) );
  AND2_X1 U454 ( .A1(n501), .A2(n521), .ZN(n380) );
  AND2_X1 U455 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U456 ( .A(KEYINPUT44), .ZN(n509) );
  INV_X1 U457 ( .A(n560), .ZN(n561) );
  INV_X1 U458 ( .A(KEYINPUT76), .ZN(n532) );
  NAND2_X1 U459 ( .A1(n421), .A2(n561), .ZN(n562) );
  INV_X1 U460 ( .A(n645), .ZN(n754) );
  INV_X1 U461 ( .A(G134), .ZN(n385) );
  INV_X1 U462 ( .A(KEYINPUT19), .ZN(n443) );
  INV_X1 U463 ( .A(KEYINPUT108), .ZN(n557) );
  BUF_X1 U464 ( .A(n565), .Z(n601) );
  INV_X1 U465 ( .A(KEYINPUT60), .ZN(n633) );
  XNOR2_X1 U466 ( .A(n626), .B(n625), .ZN(G51) );
  XOR2_X1 U467 ( .A(G137), .B(G131), .Z(n383) );
  INV_X1 U468 ( .A(KEYINPUT65), .ZN(n382) );
  XNOR2_X1 U469 ( .A(n382), .B(KEYINPUT4), .ZN(n433) );
  XNOR2_X2 U470 ( .A(n386), .B(n480), .ZN(n751) );
  XNOR2_X2 U471 ( .A(n751), .B(n387), .ZN(n403) );
  XNOR2_X1 U472 ( .A(G116), .B(G113), .ZN(n389) );
  XNOR2_X1 U473 ( .A(n390), .B(n389), .ZN(n426) );
  NOR2_X1 U474 ( .A1(G953), .A2(G237), .ZN(n468) );
  NAND2_X1 U475 ( .A1(G210), .A2(n468), .ZN(n392) );
  XNOR2_X1 U476 ( .A(KEYINPUT5), .B(G101), .ZN(n391) );
  XNOR2_X1 U477 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U478 ( .A(n426), .B(n393), .ZN(n394) );
  XNOR2_X1 U479 ( .A(n403), .B(n394), .ZN(n693) );
  INV_X1 U480 ( .A(G902), .ZN(n486) );
  NAND2_X1 U481 ( .A1(n693), .A2(n486), .ZN(n395) );
  XNOR2_X2 U482 ( .A(n395), .B(G472), .ZN(n545) );
  XNOR2_X1 U483 ( .A(n545), .B(KEYINPUT6), .ZN(n559) );
  INV_X1 U484 ( .A(n559), .ZN(n421) );
  XOR2_X1 U485 ( .A(G140), .B(KEYINPUT68), .Z(n415) );
  NAND2_X1 U486 ( .A1(G227), .A2(n756), .ZN(n396) );
  XNOR2_X1 U487 ( .A(n415), .B(n396), .ZN(n401) );
  XNOR2_X1 U488 ( .A(G101), .B(G107), .ZN(n398) );
  INV_X1 U489 ( .A(G110), .ZN(n397) );
  XNOR2_X1 U490 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U491 ( .A(G104), .B(KEYINPUT85), .ZN(n399) );
  XNOR2_X1 U492 ( .A(n400), .B(n399), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n401), .B(n427), .ZN(n402) );
  XNOR2_X1 U494 ( .A(n403), .B(n402), .ZN(n710) );
  XNOR2_X2 U495 ( .A(n404), .B(G469), .ZN(n549) );
  XNOR2_X1 U496 ( .A(G902), .B(KEYINPUT84), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n405), .B(KEYINPUT15), .ZN(n438) );
  NAND2_X1 U498 ( .A1(G234), .A2(n438), .ZN(n406) );
  XNOR2_X1 U499 ( .A(n406), .B(KEYINPUT20), .ZN(n407) );
  XNOR2_X1 U500 ( .A(KEYINPUT92), .B(n407), .ZN(n416) );
  AND2_X1 U501 ( .A1(n416), .A2(G221), .ZN(n409) );
  XNOR2_X1 U502 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n408) );
  XNOR2_X1 U503 ( .A(n409), .B(n408), .ZN(n663) );
  NAND2_X1 U504 ( .A1(G234), .A2(n756), .ZN(n410) );
  XOR2_X1 U505 ( .A(KEYINPUT8), .B(n410), .Z(n481) );
  XOR2_X1 U506 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n411) );
  XOR2_X1 U507 ( .A(G110), .B(G119), .Z(n413) );
  XNOR2_X1 U508 ( .A(G128), .B(G137), .ZN(n412) );
  XNOR2_X1 U509 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U510 ( .A(n387), .B(G125), .ZN(n434) );
  XNOR2_X1 U511 ( .A(n434), .B(KEYINPUT10), .ZN(n469) );
  XNOR2_X1 U512 ( .A(n415), .B(n469), .ZN(n750) );
  XOR2_X1 U513 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n418) );
  AND2_X1 U514 ( .A1(G217), .A2(n416), .ZN(n417) );
  XNOR2_X1 U515 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U516 ( .A1(n421), .A2(n380), .ZN(n423) );
  INV_X1 U517 ( .A(KEYINPUT33), .ZN(n422) );
  XNOR2_X1 U518 ( .A(n423), .B(n422), .ZN(n683) );
  XNOR2_X1 U519 ( .A(KEYINPUT69), .B(KEYINPUT16), .ZN(n424) );
  XNOR2_X1 U520 ( .A(n424), .B(G122), .ZN(n425) );
  XNOR2_X1 U521 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U522 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n430) );
  NAND2_X1 U523 ( .A1(n756), .A2(G224), .ZN(n429) );
  XNOR2_X1 U524 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U525 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U526 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n436), .B(n435), .ZN(n437) );
  INV_X1 U528 ( .A(n438), .ZN(n531) );
  NOR2_X1 U529 ( .A1(G237), .A2(G902), .ZN(n439) );
  XNOR2_X1 U530 ( .A(n439), .B(KEYINPUT70), .ZN(n441) );
  INV_X1 U531 ( .A(G210), .ZN(n617) );
  INV_X1 U532 ( .A(G214), .ZN(n440) );
  OR2_X1 U533 ( .A1(n441), .A2(n440), .ZN(n652) );
  INV_X1 U534 ( .A(n652), .ZN(n442) );
  NOR2_X2 U535 ( .A1(n565), .A2(n442), .ZN(n444) );
  NAND2_X1 U536 ( .A1(G234), .A2(G237), .ZN(n445) );
  XNOR2_X1 U537 ( .A(n445), .B(KEYINPUT14), .ZN(n448) );
  NAND2_X1 U538 ( .A1(n448), .A2(G902), .ZN(n446) );
  XNOR2_X1 U539 ( .A(n446), .B(KEYINPUT87), .ZN(n534) );
  NOR2_X1 U540 ( .A1(G898), .A2(n756), .ZN(n746) );
  NAND2_X1 U541 ( .A1(n534), .A2(n746), .ZN(n447) );
  XOR2_X1 U542 ( .A(KEYINPUT88), .B(n447), .Z(n451) );
  NAND2_X1 U543 ( .A1(n448), .A2(G952), .ZN(n450) );
  INV_X1 U544 ( .A(KEYINPUT86), .ZN(n449) );
  XNOR2_X1 U545 ( .A(n450), .B(n449), .ZN(n681) );
  AND2_X1 U546 ( .A1(n681), .A2(n756), .ZN(n537) );
  NOR2_X1 U547 ( .A1(n451), .A2(n537), .ZN(n452) );
  XNOR2_X1 U548 ( .A(n452), .B(KEYINPUT89), .ZN(n453) );
  NAND2_X1 U549 ( .A1(n577), .A2(n453), .ZN(n456) );
  INV_X1 U550 ( .A(KEYINPUT81), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n454), .B(KEYINPUT0), .ZN(n455) );
  INV_X1 U552 ( .A(KEYINPUT34), .ZN(n457) );
  XNOR2_X1 U553 ( .A(n458), .B(n457), .ZN(n490) );
  XOR2_X1 U554 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n460) );
  XNOR2_X1 U555 ( .A(G140), .B(KEYINPUT97), .ZN(n459) );
  XNOR2_X1 U556 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U557 ( .A(n461), .B(KEYINPUT98), .Z(n467) );
  XOR2_X1 U558 ( .A(KEYINPUT12), .B(G122), .Z(n463) );
  XNOR2_X1 U559 ( .A(G113), .B(G104), .ZN(n462) );
  XNOR2_X1 U560 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U561 ( .A(G143), .B(G131), .ZN(n464) );
  XNOR2_X1 U562 ( .A(n467), .B(n466), .ZN(n472) );
  NAND2_X1 U563 ( .A1(G214), .A2(n468), .ZN(n470) );
  XOR2_X1 U564 ( .A(n470), .B(n469), .Z(n471) );
  XNOR2_X1 U565 ( .A(n472), .B(n471), .ZN(n629) );
  NAND2_X1 U566 ( .A1(n629), .A2(n486), .ZN(n476) );
  XOR2_X1 U567 ( .A(KEYINPUT100), .B(KEYINPUT13), .Z(n474) );
  XNOR2_X1 U568 ( .A(KEYINPUT99), .B(G475), .ZN(n473) );
  XNOR2_X1 U569 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X2 U570 ( .A(n476), .B(n475), .ZN(n515) );
  XOR2_X1 U571 ( .A(KEYINPUT7), .B(G122), .Z(n478) );
  XNOR2_X1 U572 ( .A(G116), .B(G107), .ZN(n477) );
  XNOR2_X1 U573 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U574 ( .A(n480), .B(n479), .Z(n485) );
  NAND2_X1 U575 ( .A1(G217), .A2(n481), .ZN(n483) );
  XNOR2_X1 U576 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n704) );
  NAND2_X1 U579 ( .A1(n704), .A2(n486), .ZN(n488) );
  XNOR2_X1 U580 ( .A(KEYINPUT102), .B(G478), .ZN(n487) );
  XNOR2_X1 U581 ( .A(n488), .B(n487), .ZN(n516) );
  INV_X1 U582 ( .A(n516), .ZN(n494) );
  OR2_X1 U583 ( .A1(n515), .A2(n494), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n489), .B(KEYINPUT107), .ZN(n568) );
  NAND2_X1 U585 ( .A1(n490), .A2(n568), .ZN(n492) );
  XNOR2_X1 U586 ( .A(KEYINPUT71), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U587 ( .A(n492), .B(n491), .ZN(n691) );
  INV_X1 U588 ( .A(n493), .ZN(n496) );
  NAND2_X1 U589 ( .A1(n515), .A2(n494), .ZN(n655) );
  INV_X1 U590 ( .A(n663), .ZN(n495) );
  NAND2_X1 U591 ( .A1(n496), .A2(n379), .ZN(n499) );
  INV_X1 U592 ( .A(KEYINPUT66), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n497), .B(KEYINPUT22), .ZN(n498) );
  INV_X1 U594 ( .A(n501), .ZN(n667) );
  NOR2_X1 U595 ( .A1(n662), .A2(n667), .ZN(n502) );
  NAND2_X1 U596 ( .A1(n511), .A2(n502), .ZN(n503) );
  INV_X1 U597 ( .A(n504), .ZN(n507) );
  OR2_X1 U598 ( .A1(n662), .A2(n501), .ZN(n505) );
  OR2_X1 U599 ( .A1(n545), .A2(n505), .ZN(n506) );
  OR2_X1 U600 ( .A1(n507), .A2(n506), .ZN(n635) );
  AND2_X1 U601 ( .A1(n636), .A2(n635), .ZN(n508) );
  NAND2_X1 U602 ( .A1(n691), .A2(n508), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n510), .B(n509), .ZN(n526) );
  INV_X1 U604 ( .A(n511), .ZN(n512) );
  XOR2_X1 U605 ( .A(n514), .B(KEYINPUT104), .Z(n735) );
  INV_X1 U606 ( .A(n735), .ZN(n725) );
  NOR2_X2 U607 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X2 U608 ( .A(n517), .B(KEYINPUT103), .ZN(n558) );
  NAND2_X1 U609 ( .A1(n725), .A2(n558), .ZN(n518) );
  XNOR2_X1 U610 ( .A(n657), .B(KEYINPUT74), .ZN(n584) );
  NAND2_X1 U611 ( .A1(n545), .A2(n380), .ZN(n672) );
  OR2_X1 U612 ( .A1(n493), .A2(n672), .ZN(n520) );
  XOR2_X1 U613 ( .A(KEYINPUT31), .B(KEYINPUT95), .Z(n519) );
  XNOR2_X1 U614 ( .A(n520), .B(n519), .ZN(n734) );
  INV_X1 U615 ( .A(n539), .ZN(n522) );
  OR2_X1 U616 ( .A1(n545), .A2(n522), .ZN(n523) );
  NOR2_X1 U617 ( .A1(n493), .A2(n523), .ZN(n720) );
  NOR2_X1 U618 ( .A1(n734), .A2(n720), .ZN(n524) );
  OR2_X1 U619 ( .A1(n584), .A2(n524), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n381), .A2(n526), .ZN(n530) );
  XNOR2_X1 U621 ( .A(KEYINPUT78), .B(KEYINPUT45), .ZN(n528) );
  INV_X1 U622 ( .A(KEYINPUT64), .ZN(n527) );
  XNOR2_X1 U623 ( .A(n528), .B(n527), .ZN(n529) );
  NAND2_X1 U624 ( .A1(n610), .A2(n531), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n533), .B(n532), .ZN(n607) );
  NAND2_X1 U626 ( .A1(G953), .A2(n534), .ZN(n535) );
  NOR2_X1 U627 ( .A1(G900), .A2(n535), .ZN(n536) );
  NOR2_X1 U628 ( .A1(n537), .A2(n536), .ZN(n546) );
  NOR2_X1 U629 ( .A1(n546), .A2(n540), .ZN(n543) );
  NAND2_X1 U630 ( .A1(n545), .A2(n652), .ZN(n541) );
  XOR2_X1 U631 ( .A(KEYINPUT30), .B(n541), .Z(n542) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT38), .ZN(n653) );
  XNOR2_X1 U633 ( .A(n544), .B(KEYINPUT40), .ZN(n761) );
  INV_X1 U634 ( .A(n545), .ZN(n666) );
  NOR2_X1 U635 ( .A1(n546), .A2(n662), .ZN(n547) );
  NAND2_X1 U636 ( .A1(n663), .A2(n547), .ZN(n560) );
  NOR2_X1 U637 ( .A1(n666), .A2(n560), .ZN(n548) );
  XOR2_X1 U638 ( .A(KEYINPUT28), .B(n548), .Z(n551) );
  INV_X1 U639 ( .A(n549), .ZN(n550) );
  NOR2_X1 U640 ( .A1(n551), .A2(n550), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n653), .A2(n652), .ZN(n656) );
  XNOR2_X1 U642 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n552) );
  INV_X1 U643 ( .A(n684), .ZN(n554) );
  NAND2_X1 U644 ( .A1(n576), .A2(n554), .ZN(n555) );
  NOR2_X1 U645 ( .A1(n761), .A2(n760), .ZN(n556) );
  XNOR2_X1 U646 ( .A(n556), .B(KEYINPUT46), .ZN(n594) );
  INV_X1 U647 ( .A(n564), .ZN(n598) );
  XNOR2_X1 U648 ( .A(n566), .B(KEYINPUT36), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n567), .A2(n501), .ZN(n737) );
  INV_X1 U650 ( .A(n737), .ZN(n583) );
  INV_X1 U651 ( .A(n568), .ZN(n569) );
  NOR2_X1 U652 ( .A1(n569), .A2(n601), .ZN(n570) );
  NAND2_X1 U653 ( .A1(n571), .A2(n570), .ZN(n639) );
  NAND2_X1 U654 ( .A1(n657), .A2(KEYINPUT47), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n639), .A2(n572), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n573), .A2(KEYINPUT73), .ZN(n575) );
  INV_X1 U657 ( .A(KEYINPUT73), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n639), .A2(n586), .ZN(n574) );
  NAND2_X1 U659 ( .A1(n575), .A2(n574), .ZN(n581) );
  AND2_X1 U660 ( .A1(n577), .A2(n576), .ZN(n729) );
  INV_X1 U661 ( .A(n729), .ZN(n726) );
  NOR2_X1 U662 ( .A1(n726), .A2(KEYINPUT47), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n584), .A2(KEYINPUT67), .ZN(n578) );
  NAND2_X1 U664 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U665 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U666 ( .A1(n583), .A2(n582), .ZN(n592) );
  INV_X1 U667 ( .A(n584), .ZN(n585) );
  NAND2_X1 U668 ( .A1(KEYINPUT67), .A2(n585), .ZN(n589) );
  AND2_X1 U669 ( .A1(n586), .A2(n657), .ZN(n587) );
  NOR2_X1 U670 ( .A1(n726), .A2(n587), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n590), .A2(KEYINPUT47), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(n595), .ZN(n611) );
  NOR2_X1 U675 ( .A1(n597), .A2(n725), .ZN(n740) );
  INV_X1 U676 ( .A(n740), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT109), .B(n598), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n599), .A2(n667), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT43), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n638) );
  AND2_X1 U681 ( .A1(n603), .A2(n638), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n611), .A2(n604), .ZN(n606) );
  INV_X1 U683 ( .A(KEYINPUT77), .ZN(n605) );
  XNOR2_X2 U684 ( .A(n606), .B(n605), .ZN(n645) );
  NAND2_X1 U685 ( .A1(n607), .A2(n754), .ZN(n609) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n612) );
  OR2_X1 U687 ( .A1(n438), .A2(n612), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n611), .A2(n638), .ZN(n615) );
  OR2_X1 U689 ( .A1(n740), .A2(n612), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(KEYINPUT72), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  AND2_X1 U692 ( .A1(n352), .A2(n616), .ZN(n650) );
  INV_X1 U693 ( .A(n650), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n628), .A2(n627), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n619) );
  XNOR2_X1 U696 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n622), .B(n621), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n756), .A2(G952), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT83), .ZN(n713) );
  NAND2_X1 U700 ( .A1(n624), .A2(n713), .ZN(n626) );
  INV_X1 U701 ( .A(KEYINPUT56), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n707), .A2(G475), .ZN(n631) );
  XOR2_X1 U703 ( .A(KEYINPUT59), .B(n629), .Z(n630) );
  XNOR2_X1 U704 ( .A(n631), .B(n630), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n632), .A2(n713), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(G60) );
  XNOR2_X1 U707 ( .A(n635), .B(G110), .ZN(G12) );
  XNOR2_X1 U708 ( .A(n636), .B(G119), .ZN(G21) );
  XNOR2_X1 U709 ( .A(G140), .B(KEYINPUT118), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(G42) );
  XNOR2_X1 U711 ( .A(n639), .B(G143), .ZN(G45) );
  NOR2_X1 U712 ( .A1(n645), .A2(n641), .ZN(n644) );
  INV_X1 U713 ( .A(KEYINPUT75), .ZN(n642) );
  AND2_X1 U714 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  OR2_X2 U715 ( .A1(n644), .A2(n643), .ZN(n649) );
  NOR2_X1 U716 ( .A1(n642), .A2(KEYINPUT2), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n754), .A2(n646), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n690) );
  NOR2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n660) );
  NOR2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U723 ( .A(n658), .B(KEYINPUT120), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n661), .A2(n683), .ZN(n677) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U727 ( .A(n664), .B(KEYINPUT49), .ZN(n665) );
  NAND2_X1 U728 ( .A1(n666), .A2(n665), .ZN(n670) );
  XOR2_X1 U729 ( .A(KEYINPUT50), .B(n668), .Z(n669) );
  NOR2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n671), .B(KEYINPUT119), .ZN(n673) );
  NAND2_X1 U732 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U733 ( .A(KEYINPUT51), .B(n674), .ZN(n675) );
  NOR2_X1 U734 ( .A1(n675), .A2(n684), .ZN(n676) );
  NOR2_X1 U735 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U736 ( .A(n678), .B(KEYINPUT121), .Z(n680) );
  INV_X1 U737 ( .A(KEYINPUT52), .ZN(n679) );
  XNOR2_X1 U738 ( .A(n680), .B(n679), .ZN(n682) );
  NAND2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n688) );
  NOR2_X1 U740 ( .A1(n684), .A2(n683), .ZN(n686) );
  INV_X1 U741 ( .A(KEYINPUT122), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U743 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U744 ( .A(n691), .B(G122), .ZN(G24) );
  XNOR2_X1 U745 ( .A(n692), .B(G101), .ZN(G3) );
  NAND2_X1 U746 ( .A1(n707), .A2(G472), .ZN(n695) );
  XNOR2_X1 U747 ( .A(n693), .B(KEYINPUT62), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U749 ( .A1(n696), .A2(n713), .ZN(n698) );
  XNOR2_X1 U750 ( .A(KEYINPUT82), .B(KEYINPUT63), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n698), .B(n697), .ZN(G57) );
  NAND2_X1 U752 ( .A1(n350), .A2(G217), .ZN(n701) );
  XOR2_X1 U753 ( .A(KEYINPUT126), .B(n699), .Z(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  INV_X1 U755 ( .A(n713), .ZN(n705) );
  NOR2_X1 U756 ( .A1(n702), .A2(n705), .ZN(G66) );
  NAND2_X1 U757 ( .A1(n350), .A2(G478), .ZN(n703) );
  XOR2_X1 U758 ( .A(n704), .B(n703), .Z(n706) );
  NOR2_X1 U759 ( .A1(n706), .A2(n705), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n707), .A2(G469), .ZN(n712) );
  XNOR2_X1 U761 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n708) );
  XNOR2_X1 U762 ( .A(n708), .B(KEYINPUT58), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n715), .B(KEYINPUT125), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n732), .A2(n720), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n716), .B(KEYINPUT112), .ZN(n717) );
  XNOR2_X1 U769 ( .A(G104), .B(n717), .ZN(G6) );
  XOR2_X1 U770 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n719) );
  XNOR2_X1 U771 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n724) );
  XNOR2_X1 U773 ( .A(G107), .B(KEYINPUT26), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n720), .A2(n735), .ZN(n721) );
  XNOR2_X1 U775 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n724), .B(n723), .ZN(G9) );
  NOR2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U778 ( .A(G128), .B(KEYINPUT29), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(G30) );
  NAND2_X1 U780 ( .A1(n729), .A2(n732), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n730), .B(KEYINPUT116), .ZN(n731) );
  XNOR2_X1 U782 ( .A(G146), .B(n731), .ZN(G48) );
  NAND2_X1 U783 ( .A1(n732), .A2(n734), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(G113), .ZN(G15) );
  NAND2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n736), .B(G116), .ZN(G18) );
  XNOR2_X1 U787 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(G125), .B(n739), .ZN(G27) );
  XOR2_X1 U790 ( .A(G134), .B(n740), .Z(G36) );
  NAND2_X1 U791 ( .A1(n352), .A2(n756), .ZN(n744) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n741) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n741), .ZN(n742) );
  NAND2_X1 U794 ( .A1(n742), .A2(G898), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n749) );
  XOR2_X1 U796 ( .A(KEYINPUT127), .B(n745), .Z(n747) );
  NOR2_X1 U797 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n749), .B(n748), .ZN(G69) );
  XNOR2_X1 U799 ( .A(n751), .B(n750), .ZN(n755) );
  XNOR2_X1 U800 ( .A(G227), .B(n755), .ZN(n752) );
  NAND2_X1 U801 ( .A1(G900), .A2(n752), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(G953), .ZN(n759) );
  XNOR2_X1 U803 ( .A(n755), .B(n645), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n759), .A2(n758), .ZN(G72) );
  XOR2_X1 U806 ( .A(G137), .B(n760), .Z(G39) );
  XOR2_X1 U807 ( .A(G131), .B(n761), .Z(G33) );
endmodule

