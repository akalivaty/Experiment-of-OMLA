//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(G137), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XOR2_X1   g050(.A(KEYINPUT3), .B(G2104), .Z(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n467), .A2(new_n469), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n483), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n470), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n474), .B1(new_n482), .B2(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n465), .A2(new_n479), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n465), .A2(new_n466), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND3_X1  g071(.A1(new_n470), .A2(new_n483), .A3(G138), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n497), .A2(new_n498), .B1(G102), .B2(new_n472), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n463), .B2(new_n464), .ZN(new_n501));
  AND2_X1   g076(.A1(G114), .A2(G2104), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n499), .A2(KEYINPUT69), .A3(new_n503), .A4(new_n504), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT70), .B(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT71), .B(G651), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(G50), .A3(G543), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(G88), .A3(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n513), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n520), .A2(new_n527), .A3(new_n529), .ZN(G166));
  NAND4_X1  g105(.A1(new_n514), .A2(G89), .A3(new_n518), .A4(new_n526), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n514), .A2(G51), .A3(new_n518), .A4(G543), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n522), .A2(new_n524), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  AND4_X1   g113(.A1(new_n531), .A2(new_n532), .A3(new_n536), .A4(new_n538), .ZN(G168));
  NAND4_X1  g114(.A1(new_n514), .A2(G90), .A3(new_n518), .A4(new_n526), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n514), .A2(G52), .A3(new_n518), .A4(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n525), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND3_X1  g122(.A1(new_n522), .A2(new_n524), .A3(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n548), .A2(new_n552), .A3(new_n549), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(G651), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n514), .A2(G81), .A3(new_n518), .A4(new_n526), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n514), .A2(G43), .A3(new_n518), .A4(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT74), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n554), .A2(new_n559), .A3(new_n555), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND4_X1  g142(.A1(new_n514), .A2(G91), .A3(new_n518), .A4(new_n526), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n525), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n570), .A2(new_n571), .B1(G651), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n514), .A2(G53), .A3(new_n518), .A4(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G299));
  NAND4_X1  g153(.A1(new_n531), .A2(new_n532), .A3(new_n536), .A4(new_n538), .ZN(G286));
  NAND3_X1  g154(.A1(new_n520), .A2(new_n527), .A3(new_n529), .ZN(G303));
  NAND3_X1  g155(.A1(new_n519), .A2(G49), .A3(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n514), .A2(G87), .A3(new_n518), .A4(new_n526), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n526), .A2(new_n585), .A3(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT76), .B1(new_n525), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n519), .A2(new_n526), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(G305));
  INV_X1    g170(.A(new_n593), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n519), .A2(G543), .ZN(new_n597));
  AOI22_X1  g172(.A1(G85), .A2(new_n596), .B1(new_n597), .B2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n525), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(G651), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n598), .A2(new_n607), .A3(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n514), .A2(G92), .A3(new_n518), .A4(new_n526), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n514), .A2(G54), .A3(new_n518), .A4(G543), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n525), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G651), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n615), .B1(new_n614), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n613), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n610), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G299), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G860), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n622), .B1(G559), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT80), .Z(G148));
  INV_X1    g207(.A(new_n561), .ZN(new_n633));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n622), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n483), .A2(new_n472), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  OAI221_X1 g217(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n643));
  INV_X1    g218(.A(G123), .ZN(new_n644));
  INV_X1    g219(.A(G135), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n643), .B1(new_n488), .B2(new_n644), .C1(new_n645), .C2(new_n491), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT81), .B(G2438), .Z(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT15), .B(G2435), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(G14), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT82), .Z(new_n669));
  XOR2_X1   g244(.A(new_n667), .B(KEYINPUT17), .Z(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n667), .A3(new_n663), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n665), .A3(new_n663), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n685), .A2(new_n686), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n682), .A2(new_n687), .A3(new_n684), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(new_n686), .C2(new_n685), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT84), .B(G1981), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n699));
  INV_X1    g274(.A(G24), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G290), .B2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n703), .B2(new_n699), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(new_n691), .ZN(new_n705));
  OAI211_X1 g280(.A(G1986), .B(new_n701), .C1(new_n703), .C2(new_n699), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI221_X1 g282(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n708));
  INV_X1    g283(.A(G119), .ZN(new_n709));
  INV_X1    g284(.A(G131), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n708), .B1(new_n488), .B2(new_n709), .C1(new_n710), .C2(new_n491), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G23), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G288), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT33), .B(G1976), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(KEYINPUT86), .B(new_n717), .C1(G288), .C2(G16), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n721), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n722), .B1(new_n720), .B2(new_n724), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(G16), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G303), .B2(new_n716), .ZN(new_n730));
  INV_X1    g305(.A(G1971), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g307(.A(G1971), .B(new_n729), .C1(G303), .C2(new_n716), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(G305), .A2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G6), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT32), .B(G1981), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n735), .B(new_n738), .C1(new_n736), .C2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n734), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n728), .A2(new_n742), .A3(KEYINPUT34), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT34), .B1(new_n728), .B2(new_n742), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n707), .B(new_n715), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n746));
  OAI21_X1  g321(.A(KEYINPUT88), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n715), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n728), .A2(new_n742), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n728), .A2(new_n742), .A3(KEYINPUT34), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n754));
  INV_X1    g329(.A(new_n746), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n707), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n745), .A2(KEYINPUT36), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n747), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n716), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n716), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT94), .B(G1966), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n763));
  INV_X1    g338(.A(G34), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(new_n474), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n485), .A2(KEYINPUT67), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n484), .A2(new_n481), .A3(new_n470), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n770), .B(new_n771), .C1(new_n775), .C2(new_n766), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G5), .B2(G16), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n779), .A2(G5), .A3(G16), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n780), .B(new_n781), .C1(G301), .C2(new_n716), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n472), .A2(G105), .ZN(new_n787));
  INV_X1    g362(.A(G141), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n786), .B(new_n787), .C1(new_n491), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G129), .B2(new_n489), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G29), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G29), .B2(G32), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT27), .B(G1996), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n778), .B(new_n784), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n795));
  INV_X1    g370(.A(G11), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n762), .B(new_n795), .C1(KEYINPUT31), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n782), .A2(new_n783), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n766), .A2(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n766), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT29), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2090), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n797), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n716), .A2(KEYINPUT23), .A3(G20), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT23), .ZN(new_n809));
  INV_X1    g384(.A(G20), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(G16), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n811), .C1(new_n627), .C2(new_n716), .ZN(new_n812));
  INV_X1    g387(.A(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n623), .A2(new_n716), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G4), .B2(new_n716), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n817), .A2(G1348), .B1(KEYINPUT96), .B2(new_n794), .ZN(new_n818));
  NAND2_X1  g393(.A1(G115), .A2(G2104), .ZN(new_n819));
  INV_X1    g394(.A(G127), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n476), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n492), .A2(G139), .B1(new_n821), .B2(new_n479), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT25), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(KEYINPUT25), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G33), .B(new_n826), .S(G29), .Z(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G2072), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n792), .A2(new_n793), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n776), .A2(new_n777), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n814), .B(new_n818), .C1(KEYINPUT93), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n796), .A2(KEYINPUT31), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(KEYINPUT93), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n766), .A2(G26), .ZN(new_n835));
  OAI221_X1 g410(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n489), .A2(G128), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n492), .A2(G140), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n835), .B1(new_n841), .B2(G29), .ZN(new_n842));
  MUX2_X1   g417(.A(new_n835), .B(new_n842), .S(KEYINPUT28), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G2067), .ZN(new_n844));
  AND2_X1   g419(.A1(KEYINPUT30), .A2(G28), .ZN(new_n845));
  NOR2_X1   g420(.A1(KEYINPUT30), .A2(G28), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n766), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n834), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NOR4_X1   g423(.A1(new_n807), .A2(new_n832), .A3(new_n833), .A4(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n646), .A2(new_n766), .ZN(new_n850));
  NOR2_X1   g425(.A1(G16), .A2(G19), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n561), .B2(G16), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT89), .B(G1341), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n758), .A2(new_n849), .A3(new_n850), .A4(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n817), .A2(G1348), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G311));
  AND3_X1   g432(.A1(new_n758), .A2(new_n849), .A3(new_n854), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n859));
  INV_X1    g434(.A(new_n856), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n850), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT97), .B1(new_n855), .B2(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(G150));
  NAND4_X1  g438(.A1(new_n514), .A2(G55), .A3(new_n518), .A4(G543), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT98), .B(G93), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n514), .A2(new_n518), .A3(new_n526), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  INV_X1    g442(.A(G67), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n525), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G651), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n864), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n623), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT38), .ZN(new_n875));
  INV_X1    g450(.A(new_n871), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n558), .B2(new_n560), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n557), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n875), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT99), .Z(new_n884));
  OAI21_X1  g459(.A(new_n630), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n873), .B1(new_n884), .B2(new_n885), .ZN(G145));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n711), .B(new_n640), .ZN(new_n888));
  AOI22_X1  g463(.A1(G130), .A2(new_n489), .B1(new_n492), .B2(G142), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n470), .A2(G118), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT100), .Z(new_n891));
  OAI21_X1  g466(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n888), .B(new_n893), .Z(new_n894));
  AND3_X1   g469(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n841), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n826), .B(new_n790), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n894), .A3(new_n899), .ZN(new_n902));
  XNOR2_X1  g477(.A(G160), .B(new_n495), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n646), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n900), .B2(KEYINPUT101), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n898), .A2(new_n894), .A3(new_n907), .A4(new_n899), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT102), .B(new_n904), .C1(new_n906), .C2(new_n908), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n887), .B(new_n905), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(new_n871), .A2(new_n634), .ZN(new_n915));
  INV_X1    g490(.A(G305), .ZN(new_n916));
  AND2_X1   g491(.A1(G303), .A2(G288), .ZN(new_n917));
  NOR2_X1   g492(.A1(G303), .A2(G288), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n598), .A2(new_n607), .A3(new_n608), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n921));
  NAND2_X1  g496(.A1(G166), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(G303), .A2(G288), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(G305), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n919), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n928));
  NAND2_X1  g503(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n929), .B2(new_n927), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n623), .A2(new_n575), .A3(new_n577), .ZN(new_n932));
  NAND2_X1  g507(.A1(G299), .A2(new_n622), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT41), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NOR2_X1   g510(.A1(G299), .A2(new_n622), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n620), .A2(new_n621), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n937), .A2(new_n613), .B1(new_n575), .B2(new_n577), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n880), .B(new_n636), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n936), .A2(new_n938), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n941), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n931), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n915), .B1(new_n945), .B2(new_n634), .ZN(G295));
  OAI21_X1  g521(.A(new_n915), .B1(new_n945), .B2(new_n634), .ZN(G331));
  NAND2_X1  g522(.A1(new_n561), .A2(new_n871), .ZN(new_n948));
  NAND2_X1  g523(.A1(G301), .A2(KEYINPUT104), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n540), .A2(new_n541), .A3(new_n950), .A4(new_n545), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(G286), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(G168), .A2(G171), .A3(new_n950), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n954), .A3(new_n878), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n953), .B(new_n952), .C1(new_n877), .C2(new_n879), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT105), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n880), .A2(new_n958), .A3(new_n954), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n957), .A2(new_n939), .A3(new_n934), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n943), .A2(new_n955), .A3(new_n956), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n927), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n887), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n927), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT43), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n955), .A2(new_n956), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n934), .A3(new_n939), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n932), .A2(new_n933), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n957), .B2(new_n959), .ZN(new_n970));
  OAI22_X1  g545(.A1(new_n968), .A2(new_n970), .B1(new_n925), .B2(new_n926), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n887), .A4(new_n962), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT106), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  INV_X1    g554(.A(new_n970), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n927), .B1(new_n980), .B2(new_n967), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n963), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT107), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n963), .A2(new_n964), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n975), .B1(new_n984), .B2(new_n972), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(KEYINPUT43), .C1(new_n963), .C2(new_n981), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n977), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n977), .A2(KEYINPUT108), .A3(new_n979), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(G397));
  OAI211_X1 g568(.A(new_n772), .B(G40), .C1(new_n773), .C2(new_n774), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n505), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n996), .A4(new_n508), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n761), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n507), .A2(new_n996), .A3(new_n508), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(new_n994), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n777), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(G168), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G168), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1007), .B(G8), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1007), .A2(G8), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n997), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n994), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1002), .A2(new_n995), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT110), .B(G1971), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT111), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT112), .B(G2090), .Z(new_n1020));
  OR2_X1    g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1017), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G303), .A2(G8), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n591), .A2(new_n592), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT114), .B(G86), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n593), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(G1981), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(new_n1038), .C1(KEYINPUT115), .C2(KEYINPUT49), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1043));
  OAI211_X1 g618(.A(new_n1039), .B(new_n1041), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(G288), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1041), .B(new_n1048), .C1(new_n1045), .C2(G288), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1044), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1004), .B(new_n1052), .C1(new_n1002), .C2(KEYINPUT50), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1020), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1031), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1012), .A2(new_n1033), .A3(new_n1050), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(G299), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(G299), .A2(new_n1058), .A3(KEYINPUT57), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1053), .A2(new_n813), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1014), .A2(new_n1015), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  OR2_X1    g640(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(G299), .A2(new_n1058), .A3(KEYINPUT57), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n1059), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1071));
  INV_X1    g646(.A(G1996), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1014), .A2(new_n1015), .A3(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n994), .B2(new_n997), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n633), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1076), .A2(KEYINPUT121), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(KEYINPUT121), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n633), .B(new_n1079), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1067), .B(new_n1071), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n994), .A2(G2067), .A3(new_n997), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1083), .B(new_n1084), .C1(new_n1019), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n623), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1019), .B2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(KEYINPUT123), .A3(new_n622), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1088), .A2(new_n1091), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1082), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1069), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1089), .A2(new_n622), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1065), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1057), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1022), .B2(G2078), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n772), .A2(G40), .A3(new_n480), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n997), .A2(new_n995), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT126), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1099), .A2(G2078), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1103), .A2(new_n1104), .A3(new_n1110), .A4(new_n1105), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1019), .A2(KEYINPUT124), .A3(new_n783), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT124), .B1(new_n1019), .B2(new_n783), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1100), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1100), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1019), .A2(new_n783), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n998), .A2(new_n999), .A3(new_n1109), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(G171), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT54), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1115), .A2(G171), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1100), .A2(G301), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT54), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(KEYINPUT127), .A3(KEYINPUT54), .A4(new_n1124), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1098), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1033), .A2(new_n1050), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1026), .A2(G8), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1031), .ZN(new_n1135));
  AOI211_X1 g710(.A(new_n1040), .B(G286), .C1(new_n1001), .C2(new_n1006), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1131), .A2(new_n1132), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1026), .A2(G8), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT63), .B1(new_n1138), .B2(new_n1032), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1033), .A2(new_n1050), .A3(new_n1136), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1033), .A2(new_n1050), .A3(new_n1056), .A4(new_n1136), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1133), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1142), .B2(new_n1133), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1137), .B(new_n1141), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1131), .A2(new_n1056), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1121), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1138), .A2(new_n1032), .A3(new_n1050), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1044), .A2(new_n1045), .A3(new_n921), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1034), .B(KEYINPUT116), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1041), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1152), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1130), .A2(new_n1146), .A3(new_n1151), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1104), .A2(new_n994), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT109), .Z(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n841), .B(G2067), .Z(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1072), .B2(new_n790), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1161), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(G1996), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1163), .A2(new_n1165), .B1(new_n790), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n711), .B(new_n714), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(G290), .B(G1986), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1161), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1160), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1162), .B1(new_n790), .B2(new_n1164), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1167), .B(KEYINPUT46), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT47), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n711), .A2(new_n713), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1168), .A2(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n841), .A2(G2067), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1162), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1166), .A2(G290), .A3(G1986), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT48), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1170), .A2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1177), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1173), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g761(.A1(new_n913), .A2(G319), .ZN(new_n1188));
  NOR2_X1   g762(.A1(G229), .A2(G401), .ZN(new_n1189));
  NAND4_X1  g763(.A1(new_n1188), .A2(new_n677), .A3(new_n974), .A4(new_n1189), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


