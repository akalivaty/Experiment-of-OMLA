//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT84), .B(G224), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n195), .B1(new_n193), .B2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n203), .A2(new_n195), .A3(G128), .A4(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(G125), .B1(new_n198), .B2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n194), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n204), .B1(new_n193), .B2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n211), .A2(new_n213), .A3(G125), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n189), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n194), .A2(new_n210), .B1(new_n212), .B2(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n197), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n200), .A2(new_n202), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n191), .B1(new_n219), .B2(new_n190), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n206), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G125), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n189), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(G116), .A2(G119), .ZN(new_n227));
  NOR2_X1   g041(.A1(G116), .A2(G119), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n229), .B(new_n230), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT75), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G104), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n237), .A3(G107), .ZN(new_n238));
  AOI21_X1  g052(.A(G107), .B1(new_n235), .B2(new_n237), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n242), .A3(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT76), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT76), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(new_n240), .A3(new_n242), .A4(G104), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n233), .B(G101), .C1(new_n241), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G101), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n235), .A2(new_n237), .A3(G107), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n235), .A2(new_n237), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n242), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(new_n246), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n249), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT75), .B(G104), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT3), .B1(new_n256), .B2(G107), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT77), .B(G101), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n254), .A3(new_n258), .A4(new_n238), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT4), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n232), .B(new_n248), .C1(new_n255), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G119), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT80), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT81), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n264), .A2(KEYINPUT80), .ZN(new_n271));
  OAI22_X1  g085(.A1(new_n270), .A2(new_n271), .B1(new_n228), .B2(new_n227), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n263), .A2(new_n265), .A3(new_n267), .A4(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n269), .A2(G113), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G113), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n268), .B2(KEYINPUT81), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n279), .A2(KEYINPUT82), .A3(new_n272), .A4(new_n274), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n229), .A2(new_n230), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n242), .A2(G104), .ZN(new_n283));
  OAI21_X1  g097(.A(G101), .B1(new_n239), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n259), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(G110), .B(G122), .Z(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n261), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT6), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n261), .A2(new_n286), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n288), .A2(KEYINPUT83), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(KEYINPUT6), .A3(new_n292), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n226), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n224), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n215), .A2(new_n225), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n287), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n259), .A2(new_n284), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n279), .A2(new_n274), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n229), .A2(new_n264), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n282), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n303), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n281), .A2(new_n282), .A3(new_n304), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n217), .A2(new_n223), .A3(new_n299), .A4(new_n224), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n301), .A2(new_n289), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n296), .A2(new_n298), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n226), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n289), .A2(KEYINPUT6), .B1(new_n291), .B2(new_n292), .ZN(new_n318));
  INV_X1    g132(.A(new_n295), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n313), .A2(new_n314), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n297), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n187), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(G143), .A3(G214), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(G143), .B1(new_n324), .B2(G214), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n327), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n325), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n222), .A2(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n338), .B1(new_n341), .B2(new_n336), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(G146), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT88), .A4(new_n332), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n329), .A2(new_n325), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT17), .A3(G131), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n335), .A2(new_n343), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n193), .A2(new_n339), .A3(new_n340), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(G146), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT18), .A2(G131), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n345), .A2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT87), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n234), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n347), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT89), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n347), .A2(new_n360), .A3(new_n354), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(G146), .B(new_n338), .C1(new_n341), .C2(new_n336), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n341), .B(KEYINPUT19), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT86), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT86), .B1(new_n328), .B2(new_n331), .ZN(new_n366));
  OAI221_X1 g180(.A(new_n363), .B1(new_n219), .B2(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n354), .ZN(new_n368));
  INV_X1    g182(.A(new_n357), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n372));
  NOR2_X1   g186(.A1(G475), .A2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n359), .A2(new_n361), .B1(new_n369), .B2(new_n368), .ZN(new_n375));
  INV_X1    g189(.A(new_n373), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n357), .B1(new_n347), .B2(new_n354), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n359), .B2(new_n361), .ZN(new_n380));
  OAI21_X1  g194(.A(G475), .B1(new_n380), .B2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G478), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT15), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  INV_X1    g199(.A(G217), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n385), .A2(new_n386), .A3(G953), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n197), .A2(G143), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n190), .B2(G128), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n197), .A2(KEYINPUT91), .A3(G143), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT65), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G134), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G116), .B(G122), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(new_n242), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G116), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n262), .A2(G122), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G107), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n400), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT92), .ZN(new_n409));
  OR2_X1    g223(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(new_n389), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n409), .A3(new_n389), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n391), .A2(new_n392), .ZN(new_n416));
  INV_X1    g230(.A(new_n389), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n410), .A3(new_n411), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n408), .B1(new_n419), .B2(G134), .ZN(new_n420));
  INV_X1    g234(.A(new_n407), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n423));
  OAI21_X1  g237(.A(G107), .B1(new_n405), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n393), .A2(new_n399), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n400), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n388), .B1(new_n420), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n415), .A2(new_n418), .A3(new_n416), .ZN(new_n430));
  OAI21_X1  g244(.A(G134), .B1(new_n430), .B2(new_n413), .ZN(new_n431));
  INV_X1    g245(.A(new_n408), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n400), .ZN(new_n434));
  OAI221_X1 g248(.A(new_n421), .B1(new_n422), .B2(new_n424), .C1(new_n434), .C2(new_n426), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n435), .A3(new_n387), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT93), .B1(new_n437), .B2(new_n314), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n439), .B(G902), .C1(new_n429), .C2(new_n436), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n384), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT94), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n437), .B(new_n314), .C1(KEYINPUT15), .C2(new_n383), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(new_n384), .C1(new_n438), .C2(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(G234), .A2(G237), .ZN(new_n446));
  INV_X1    g260(.A(G953), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n446), .A2(G952), .A3(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT21), .B(G898), .Z(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT95), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n446), .A2(G902), .A3(G953), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n442), .A2(new_n443), .A3(new_n445), .A4(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n382), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT96), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT96), .B1(new_n382), .B2(new_n455), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n323), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G119), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G128), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(G128), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n462), .B(new_n463), .C1(new_n464), .C2(KEYINPUT23), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G110), .ZN(new_n466));
  OR3_X1    g280(.A1(new_n461), .A2(KEYINPUT71), .A3(G128), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT71), .B1(new_n461), .B2(G128), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n462), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT24), .B(G110), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n343), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(G110), .B2(new_n465), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n363), .A3(new_n348), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n447), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT22), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(G137), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n475), .A3(new_n479), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT73), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT73), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n386), .B1(G234), .B2(new_n314), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n487), .A2(G902), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n314), .A3(new_n482), .ZN(new_n491));
  NOR2_X1   g305(.A1(KEYINPUT72), .A2(KEYINPUT25), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n488), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n496), .A3(KEYINPUT74), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT74), .ZN(new_n498));
  INV_X1    g312(.A(new_n488), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n493), .B2(new_n494), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n489), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G137), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT11), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n395), .A2(new_n397), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(KEYINPUT11), .A3(G134), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G137), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n395), .A2(new_n397), .A3(new_n504), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n511), .A2(new_n330), .A3(new_n506), .A4(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(KEYINPUT66), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(G131), .C1(new_n505), .C2(new_n509), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n216), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n330), .B1(G134), .B2(G137), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n398), .B2(G137), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n221), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n519), .A3(new_n231), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n231), .B1(new_n516), .B2(new_n519), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n522), .B1(new_n527), .B2(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n519), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n232), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n520), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n528), .B1(new_n531), .B2(KEYINPUT68), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n324), .A2(G210), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n533), .B(KEYINPUT27), .Z(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT26), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n249), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n526), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT70), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n526), .A2(new_n532), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n516), .A2(new_n519), .A3(KEYINPUT30), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n232), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n536), .B1(new_n544), .B2(new_n520), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT29), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n538), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n531), .A2(KEYINPUT28), .ZN(new_n548));
  AND4_X1   g362(.A1(KEYINPUT29), .A2(new_n526), .A3(new_n536), .A4(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(G902), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(G472), .A2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n525), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n530), .A2(new_n555), .A3(new_n520), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT28), .B1(new_n530), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n523), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n536), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n544), .A2(new_n520), .A3(new_n536), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n558), .A2(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n544), .A2(new_n520), .A3(new_n536), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT67), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n544), .A2(new_n536), .A3(KEYINPUT67), .A4(new_n520), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(KEYINPUT31), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n553), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n551), .A2(G472), .B1(new_n568), .B2(KEYINPUT32), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n502), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n314), .ZN(new_n575));
  XNOR2_X1  g389(.A(G110), .B(G140), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n447), .A2(G227), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n513), .A2(new_n515), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n304), .A2(new_n198), .A3(new_n206), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n197), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n206), .B1(new_n212), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n259), .A3(new_n284), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n255), .A2(new_n260), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n248), .A2(new_n216), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT78), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n248), .A2(new_n216), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  OAI21_X1  g406(.A(G101), .B1(new_n241), .B2(new_n247), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n259), .A4(new_n284), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AND4_X1   g415(.A1(KEYINPUT79), .A2(new_n596), .A3(new_n579), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n590), .B2(new_n595), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT79), .B1(new_n603), .B2(new_n579), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n587), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n588), .A2(KEYINPUT78), .A3(new_n589), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n592), .B1(new_n591), .B2(new_n594), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n579), .B(new_n601), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n603), .A2(KEYINPUT79), .A3(new_n579), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n578), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n603), .A2(new_n579), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n578), .A2(new_n605), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n575), .B1(new_n614), .B2(G469), .ZN(new_n615));
  INV_X1    g429(.A(new_n578), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n587), .B(new_n616), .C1(new_n602), .C2(new_n604), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n603), .A2(new_n579), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n610), .B2(new_n611), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n616), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n574), .A3(new_n314), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n573), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n460), .A2(new_n571), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(new_n258), .Z(G3));
  OAI21_X1  g438(.A(new_n383), .B1(new_n438), .B2(new_n440), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n437), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n429), .A2(new_n436), .A3(KEYINPUT33), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n314), .A2(G478), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n382), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n323), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n298), .B1(new_n296), .B2(new_n315), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n320), .A2(new_n321), .A3(new_n297), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(KEYINPUT97), .A3(new_n187), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n453), .B(new_n632), .C1(new_n634), .C2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n568), .ZN(new_n641));
  INV_X1    g455(.A(G472), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n562), .B2(new_n567), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n502), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n622), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  AOI21_X1  g463(.A(KEYINPUT97), .B1(new_n637), .B2(new_n187), .ZN(new_n650));
  INV_X1    g464(.A(new_n187), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n633), .B(new_n651), .C1(new_n635), .C2(new_n636), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n378), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n381), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(KEYINPUT99), .B(G475), .C1(new_n380), .C2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n374), .A2(new_n377), .A3(KEYINPUT98), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n655), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n653), .A2(new_n453), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n646), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT35), .B(G107), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  XNOR2_X1  g481(.A(new_n476), .B(KEYINPUT100), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n488), .A2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n496), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n496), .A3(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n644), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n460), .A2(new_n679), .A3(new_n622), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NAND2_X1  g496(.A1(new_n551), .A2(G472), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n570), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n676), .A2(new_n677), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n622), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n448), .B1(new_n452), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n662), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n634), .A2(new_n638), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NAND2_X1  g510(.A1(new_n565), .A2(new_n566), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n559), .B2(new_n531), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n570), .A2(new_n684), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n700), .A2(new_n496), .A3(new_n673), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n316), .A2(new_n322), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(KEYINPUT38), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(KEYINPUT38), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n382), .A2(new_n660), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n187), .A2(new_n701), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n690), .B(KEYINPUT39), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n622), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n622), .A2(KEYINPUT102), .A3(new_n708), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(KEYINPUT40), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT40), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n707), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  NOR2_X1   g530(.A1(new_n632), .A2(new_n690), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n692), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n688), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  OAI21_X1  g535(.A(new_n613), .B1(new_n602), .B2(new_n604), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n722), .A2(new_n578), .B1(new_n612), .B2(new_n587), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n572), .A3(new_n621), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n571), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n640), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT41), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n278), .ZN(G15));
  NOR2_X1   g544(.A1(new_n664), .A2(new_n727), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n262), .ZN(G18));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n725), .B2(new_n653), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n722), .A2(new_n578), .ZN(new_n735));
  AOI211_X1 g549(.A(G469), .B(G902), .C1(new_n735), .C2(new_n617), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n574), .B1(new_n620), .B2(new_n314), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n692), .A3(KEYINPUT103), .A4(new_n572), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n458), .A2(new_n459), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n685), .A3(new_n686), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  NAND2_X1  g558(.A1(new_n692), .A2(new_n706), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n724), .A2(new_n572), .A3(new_n621), .A4(new_n454), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n526), .A2(new_n548), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n559), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n567), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n560), .A2(new_n561), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n567), .A2(new_n749), .A3(KEYINPUT105), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n552), .B(KEYINPUT104), .Z(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n489), .A2(new_n500), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n562), .A2(new_n567), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n314), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G472), .ZN(new_n761));
  AND4_X1   g575(.A1(KEYINPUT106), .A2(new_n757), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n642), .B1(new_n759), .B2(new_n314), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n755), .B2(new_n756), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT106), .B1(new_n764), .B2(new_n758), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n747), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n674), .A3(new_n717), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n734), .B2(new_n739), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n222), .ZN(G27));
  NAND2_X1  g584(.A1(new_n615), .A2(new_n621), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n637), .A2(new_n651), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n771), .A2(new_n572), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n571), .A4(new_n717), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n497), .A2(new_n501), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n685), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n771), .A2(new_n717), .A3(new_n572), .A4(new_n772), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT107), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n568), .A2(new_n782), .A3(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n568), .B2(KEYINPUT32), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n569), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n758), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n780), .A3(new_n778), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NAND3_X1  g604(.A1(new_n773), .A2(new_n571), .A3(new_n691), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  OAI211_X1 g606(.A(new_n613), .B(new_n616), .C1(new_n602), .C2(new_n604), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n586), .B1(new_n610), .B2(new_n611), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n616), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n574), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n614), .A2(KEYINPUT45), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n575), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n575), .B1(new_n797), .B2(new_n798), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT46), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n621), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n378), .A2(new_n631), .A3(new_n381), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n644), .A3(new_n674), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n806), .A2(new_n572), .A3(new_n708), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n809), .A2(new_n644), .A3(KEYINPUT44), .A4(new_n674), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n772), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(KEYINPUT109), .A3(new_n772), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n503), .ZN(G39));
  OAI21_X1  g634(.A(new_n621), .B1(new_n804), .B2(KEYINPUT46), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n802), .B(new_n575), .C1(new_n797), .C2(new_n798), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n572), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT47), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n717), .A2(new_n502), .A3(new_n772), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT110), .A3(new_n570), .A4(new_n569), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n717), .A2(new_n502), .A3(new_n772), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(new_n685), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT47), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(new_n572), .C1(new_n821), .C2(new_n822), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT111), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n824), .A2(new_n830), .A3(new_n835), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  XNOR2_X1  g652(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n690), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n445), .A2(new_n442), .A3(new_n443), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n187), .A3(new_n702), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n655), .A2(new_n661), .A3(new_n659), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT113), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n655), .A2(new_n661), .A3(new_n659), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n772), .A4(new_n842), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n685), .A2(new_n776), .A3(new_n691), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n622), .A2(new_n772), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n687), .A2(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n778), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n764), .A2(new_n674), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n764), .A2(new_n674), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT114), .B1(new_n778), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n852), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n789), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n740), .A2(new_n717), .A3(new_n854), .ZN(new_n861));
  INV_X1    g675(.A(new_n745), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n701), .A2(new_n622), .A3(new_n841), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n678), .B1(new_n569), .B2(new_n570), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n622), .B(new_n864), .C1(new_n694), .C2(new_n719), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n687), .B1(new_n693), .B2(new_n718), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n769), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n863), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n860), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n571), .B(new_n726), .C1(new_n663), .C2(new_n639), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n743), .A2(new_n766), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n743), .A2(new_n766), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n660), .A2(new_n381), .A3(new_n378), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n632), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n323), .A2(new_n453), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n645), .A2(new_n622), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n623), .A2(new_n680), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n877), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n840), .B1(new_n872), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n868), .A2(new_n871), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n571), .A2(new_n622), .A3(new_n717), .A4(new_n772), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT42), .B1(new_n888), .B2(KEYINPUT107), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n787), .B1(new_n889), .B2(new_n775), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n687), .A2(new_n849), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n855), .B1(new_n853), .B2(new_n854), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n778), .A2(new_n857), .A3(KEYINPUT114), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n891), .B(new_n791), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n874), .A2(new_n882), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n887), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n886), .A2(KEYINPUT54), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n762), .A2(new_n765), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n809), .A2(new_n448), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n772), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n824), .A2(new_n832), .B1(new_n573), .B2(new_n738), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n448), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n700), .A2(new_n502), .A3(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n725), .A2(new_n651), .A3(new_n637), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n382), .A2(new_n631), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n902), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n857), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n725), .A2(new_n705), .A3(new_n187), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n902), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT50), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n901), .A2(KEYINPUT50), .A3(new_n902), .A4(new_n917), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n921), .ZN(new_n925));
  INV_X1    g739(.A(new_n916), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n925), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n908), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT117), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n904), .B2(new_n905), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n922), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n904), .A2(new_n929), .A3(new_n905), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n907), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n912), .A2(new_n382), .A3(new_n631), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(G952), .A3(new_n447), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n915), .A2(new_n786), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT48), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n935), .B(new_n937), .C1(new_n740), .C2(new_n903), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n928), .A2(new_n933), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n882), .B1(new_n874), .B2(KEYINPUT112), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n887), .A2(new_n877), .A3(new_n940), .A4(new_n895), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT115), .B1(new_n941), .B2(new_n896), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n872), .A2(new_n885), .A3(new_n840), .ZN(new_n943));
  INV_X1    g757(.A(new_n941), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(KEYINPUT53), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(KEYINPUT115), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n900), .B(new_n939), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  OR2_X1    g762(.A1(G952), .A2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n758), .A2(new_n572), .A3(new_n187), .ZN(new_n951));
  NOR4_X1   g765(.A1(new_n700), .A2(new_n705), .A3(new_n807), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n738), .B(KEYINPUT49), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(G75));
  AOI22_X1  g769(.A1(new_n941), .A2(new_n839), .B1(new_n872), .B2(new_n897), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n314), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(G210), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT56), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n294), .A2(new_n295), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT119), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n317), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n958), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n958), .B2(new_n959), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n447), .A2(G952), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G51));
  XNOR2_X1  g781(.A(new_n575), .B(KEYINPUT57), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n956), .A2(new_n947), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n899), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n620), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n957), .A2(new_n798), .A3(new_n797), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(G54));
  NAND2_X1  g787(.A1(KEYINPUT58), .A2(G475), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT120), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n957), .A2(new_n371), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n371), .B1(new_n957), .B2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n966), .ZN(G60));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT59), .Z(new_n980));
  NOR2_X1   g794(.A1(new_n629), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n969), .B2(new_n899), .ZN(new_n982));
  INV_X1    g796(.A(new_n966), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n980), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n941), .A2(new_n839), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT53), .B1(new_n872), .B2(new_n885), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT115), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n942), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n947), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n990), .B2(new_n899), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n984), .B1(new_n991), .B2(new_n629), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n886), .B2(new_n898), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n966), .B1(new_n996), .B2(new_n487), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n941), .A2(new_n839), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n872), .A2(new_n897), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT121), .B1(new_n1000), .B2(new_n671), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT121), .ZN(new_n1002));
  INV_X1    g816(.A(new_n671), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n956), .A2(new_n1002), .A3(new_n1003), .A4(new_n994), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n997), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(KEYINPUT61), .B(new_n997), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(G66));
  OAI21_X1  g823(.A(G953), .B1(new_n451), .B2(new_n188), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n884), .A2(KEYINPUT122), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT122), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n940), .A2(new_n1012), .A3(new_n877), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n961), .B1(G898), .B2(new_n447), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G69));
  AOI21_X1  g831(.A(new_n819), .B1(new_n834), .B2(new_n836), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n786), .A2(new_n745), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1019), .A2(new_n806), .A3(new_n572), .A4(new_n708), .ZN(new_n1020));
  AND4_X1   g834(.A1(new_n789), .A2(new_n791), .A3(new_n870), .A4(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1018), .A2(new_n447), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n542), .A2(new_n543), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n364), .B(KEYINPUT123), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(G900), .B2(G953), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT125), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n447), .B1(G227), .B2(G900), .ZN(new_n1028));
  AOI22_X1  g842(.A1(new_n1022), .A2(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n879), .A2(new_n772), .ZN(new_n1030));
  AND4_X1   g844(.A1(new_n571), .A2(new_n711), .A3(new_n712), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n715), .A2(new_n870), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT62), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n715), .A2(KEYINPUT62), .A3(new_n870), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(G953), .B1(new_n1036), .B2(new_n1018), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1025), .B(KEYINPUT124), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1029), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1028), .A2(new_n1027), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1040), .B(new_n1041), .Z(G72));
  NAND3_X1  g856(.A1(new_n1014), .A2(new_n1018), .A3(new_n1036), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  AND2_X1   g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n544), .A2(new_n520), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n536), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1045), .B1(new_n697), .B2(new_n545), .ZN(new_n1049));
  OAI22_X1  g863(.A1(new_n1046), .A2(new_n1048), .B1(new_n946), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1011), .A2(new_n1013), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT126), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n1051), .A2(new_n1052), .A3(new_n1045), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1052), .B1(new_n1051), .B2(new_n1045), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1047), .A2(new_n536), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1055), .ZN(new_n1056));
  NOR3_X1   g870(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g871(.A(KEYINPUT127), .B1(new_n1057), .B2(new_n966), .ZN(new_n1058));
  INV_X1    g872(.A(KEYINPUT127), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n1051), .A2(new_n1045), .ZN(new_n1060));
  OAI21_X1  g874(.A(new_n1055), .B1(new_n1060), .B2(new_n1052), .ZN(new_n1061));
  OAI211_X1 g875(.A(new_n1059), .B(new_n983), .C1(new_n1061), .C2(new_n1053), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1050), .B1(new_n1058), .B2(new_n1062), .ZN(G57));
endmodule


