//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT67), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT69), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  OR4_X1    g028(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n465), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n467), .A2(new_n468), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n477), .A2(new_n465), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(new_n487), .A2(G126), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n465), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n470), .A2(KEYINPUT4), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n470), .B2(new_n496), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT72), .B(G651), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g079(.A(new_n504), .B(KEYINPUT74), .Z(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n500), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(G88), .ZN(new_n512));
  AOI22_X1  g087(.A1(G50), .A2(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n505), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT75), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n500), .A2(new_n518), .A3(G63), .A4(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT72), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT72), .A2(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT6), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n506), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(G89), .A3(new_n500), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT76), .B1(new_n507), .B2(new_n508), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n525), .A2(new_n531), .A3(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n529), .B1(G51), .B2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n530), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n510), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(new_n502), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n525), .A2(G90), .A3(new_n500), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n536), .A2(new_n542), .A3(KEYINPUT77), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n531), .B1(new_n525), .B2(G543), .ZN(new_n545));
  AOI211_X1 g120(.A(KEYINPUT76), .B(new_n508), .C1(new_n523), .C2(new_n524), .ZN(new_n546));
  OAI21_X1  g121(.A(G52), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n511), .A2(G90), .B1(new_n539), .B2(new_n502), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n543), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n530), .B2(new_n532), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n525), .A2(new_n500), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n554), .A2(new_n555), .B1(new_n503), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n564));
  OR2_X1    g139(.A1(KEYINPUT72), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(KEYINPUT72), .A2(G651), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n567), .C2(new_n506), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT78), .B1(new_n507), .B2(new_n510), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n525), .A2(new_n571), .A3(new_n500), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(G91), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n500), .B2(G65), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  INV_X1    g151(.A(G651), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n569), .A2(new_n573), .A3(new_n580), .ZN(G299));
  OAI21_X1  g156(.A(G51), .B1(new_n545), .B2(new_n546), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n582), .A2(new_n526), .A3(new_n520), .A4(new_n528), .ZN(G286));
  NAND3_X1  g158(.A1(new_n570), .A2(G87), .A3(new_n572), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n570), .A2(KEYINPUT80), .A3(G87), .A4(new_n572), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n525), .A2(G49), .A3(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n510), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n509), .A2(G48), .B1(new_n596), .B2(new_n502), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n570), .A2(G86), .A3(new_n572), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n533), .A2(G47), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n510), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n511), .A2(G85), .B1(new_n603), .B2(new_n502), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G290));
  NAND3_X1  g180(.A1(new_n570), .A2(G92), .A3(new_n572), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .A4(new_n572), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n510), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n533), .A2(G54), .B1(G651), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n615), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g191(.A(new_n615), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(new_n615), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n482), .A2(G135), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G2105), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n487), .B2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n636), .A3(new_n633), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND4_X1  g219(.A1(new_n635), .A2(new_n637), .A3(new_n643), .A4(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT82), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n652), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(G14), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT83), .Z(G401));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n642), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n636), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT20), .Z(new_n683));
  AOI211_X1 g258(.A(new_n681), .B(new_n683), .C1(new_n676), .C2(new_n680), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT84), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  NOR2_X1   g268(.A1(G5), .A2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT92), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(G301), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1961), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT24), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n701), .B2(G34), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G160), .B2(G29), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n700), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n482), .A2(G141), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n487), .A2(G129), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT26), .Z(new_n709));
  NAND3_X1  g284(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n706), .A2(new_n707), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n699), .B1(G2084), .B2(new_n704), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT25), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  INV_X1    g294(.A(G139), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n718), .B1(new_n465), .B2(new_n719), .C1(new_n481), .C2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(G33), .B(new_n721), .S(G29), .Z(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G2072), .Z(new_n723));
  AOI22_X1  g298(.A1(new_n712), .A2(new_n713), .B1(G2084), .B2(new_n704), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT90), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n700), .A2(G26), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n482), .A2(G140), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT89), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G128), .B2(new_n487), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2067), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G19), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n558), .B2(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G1341), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(G1341), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n700), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n700), .ZN(new_n742));
  INV_X1    g317(.A(G2078), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n736), .A2(new_n739), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n726), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n747));
  NOR2_X1   g322(.A1(G4), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n622), .B2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT88), .B(G1348), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AND4_X1   g326(.A1(new_n715), .A2(new_n746), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n696), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n696), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT91), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT30), .B(G28), .ZN(new_n758));
  OR2_X1    g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n758), .A2(new_n700), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n761), .B1(new_n700), .B2(new_n634), .C1(new_n697), .C2(new_n698), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n700), .A2(G35), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT95), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n489), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2090), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n696), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n619), .B2(new_n696), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT98), .Z(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(G1956), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(G1956), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n772), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n764), .B2(new_n763), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n752), .A2(new_n765), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G23), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT85), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT86), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n588), .B2(new_n592), .ZN(new_n785));
  AOI211_X1 g360(.A(KEYINPUT86), .B(new_n591), .C1(new_n586), .C2(new_n587), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n783), .B1(new_n787), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT87), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n696), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n696), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n696), .A2(G6), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G305), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n797), .A2(new_n799), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n795), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n791), .A2(new_n792), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  INV_X1    g380(.A(G290), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n696), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n696), .B2(G24), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(G1986), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(G1986), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n487), .A2(G119), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n465), .A2(G107), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(G131), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n812), .B1(new_n813), .B2(new_n814), .C1(new_n481), .C2(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G25), .B(new_n816), .S(G29), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n810), .A2(new_n811), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n804), .A2(new_n805), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n781), .B1(new_n823), .B2(new_n824), .ZN(G311));
  XNOR2_X1  g400(.A(new_n822), .B(KEYINPUT36), .ZN(new_n826));
  INV_X1    g401(.A(new_n781), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  NOR2_X1   g403(.A1(new_n615), .A2(new_n623), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n530), .B2(new_n532), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n554), .A2(new_n833), .B1(new_n503), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n558), .A2(new_n836), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n557), .A2(new_n553), .B1(new_n832), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n830), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n836), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n487), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n465), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(G142), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n848), .B1(new_n849), .B2(new_n850), .C1(new_n481), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n639), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n734), .B(new_n721), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n711), .B(G164), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n816), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G160), .B(KEYINPUT99), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n489), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n634), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n859), .B2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g441(.A(G303), .B(G305), .Z(new_n867));
  NAND2_X1  g442(.A1(G288), .A2(KEYINPUT86), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n588), .A2(new_n784), .A3(new_n592), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n806), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(G290), .B1(new_n785), .B2(new_n786), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT102), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT102), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n867), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n867), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n610), .A2(G299), .A3(new_n614), .ZN(new_n881));
  AOI21_X1  g456(.A(G299), .B1(new_n610), .B2(new_n614), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n615), .A2(new_n619), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n610), .A2(G299), .A3(new_n614), .ZN(new_n885));
  XOR2_X1   g460(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n885), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n625), .B(new_n839), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n889), .B(new_n890), .S(new_n891), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n879), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n879), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G868), .B2(new_n836), .ZN(G295));
  OAI21_X1  g472(.A(new_n896), .B1(G868), .B2(new_n836), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT77), .B1(new_n536), .B2(new_n542), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n547), .A2(new_n548), .A3(new_n544), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n900), .A2(G286), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G286), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n839), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(G168), .B1(new_n543), .B2(new_n549), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(G286), .A3(new_n901), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n905), .A2(new_n838), .A3(new_n837), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n907), .A3(new_n890), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n889), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n904), .A2(new_n907), .A3(new_n890), .A4(KEYINPUT103), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n878), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n890), .A2(new_n887), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n884), .A2(new_n880), .A3(new_n885), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n911), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n904), .A2(new_n907), .A3(new_n890), .A4(KEYINPUT105), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n874), .A3(new_n877), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n915), .A2(new_n916), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n916), .B1(new_n915), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n904), .A2(new_n907), .A3(new_n890), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n928), .A2(KEYINPUT103), .B1(new_n889), .B2(new_n911), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n806), .B1(new_n868), .B2(new_n869), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n785), .A2(new_n786), .A3(G290), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n875), .B1(new_n933), .B2(new_n876), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n872), .A2(new_n867), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n910), .B(new_n929), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n874), .A3(new_n877), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n899), .B1(new_n927), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n936), .A2(new_n937), .A3(new_n924), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n944), .A2(KEYINPUT104), .B1(new_n945), .B2(new_n941), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n915), .B2(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT44), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT107), .B1(new_n943), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n915), .A2(new_n924), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n915), .A2(new_n916), .A3(new_n924), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n941), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n942), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n947), .A2(new_n948), .B1(new_n952), .B2(KEYINPUT43), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n944), .A2(KEYINPUT104), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n899), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n951), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G164), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G160), .A2(G40), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT109), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(G164), .B2(G1384), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND3_X1  g548(.A1(G160), .A2(new_n973), .A3(G40), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(new_n970), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n756), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n970), .A2(new_n974), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n980));
  NOR2_X1   g555(.A1(G164), .A2(G1384), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT116), .B(G2084), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n979), .A2(new_n980), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(KEYINPUT115), .A3(new_n756), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n978), .A2(new_n985), .A3(G168), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G8), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n978), .A2(new_n986), .A3(new_n985), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G286), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(G8), .A3(new_n987), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n993), .B2(KEYINPUT51), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT62), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT124), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n983), .A2(new_n970), .A3(new_n980), .A4(new_n974), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n977), .A2(new_n976), .B1(new_n998), .B2(new_n984), .ZN(new_n999));
  AOI21_X1  g574(.A(G168), .B1(new_n999), .B2(new_n986), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n987), .A2(G8), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT51), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n989), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT124), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT62), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n994), .A2(new_n995), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT55), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n966), .B1(G164), .B2(G1384), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n970), .A3(new_n1012), .A4(new_n974), .ZN(new_n1013));
  INV_X1    g588(.A(G1971), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(G2090), .B2(new_n997), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n981), .A2(new_n970), .A3(new_n974), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT113), .B(G86), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n511), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n597), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G1981), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G305), .B2(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1021), .A2(new_n1029), .A3(KEYINPUT114), .A4(new_n1028), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n787), .A2(G1976), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1021), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1021), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1034), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1008), .ZN(new_n1042));
  INV_X1    g617(.A(new_n982), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(G164), .B2(G1384), .ZN(new_n1044));
  OR3_X1    g619(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n979), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1046), .A2(G2090), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1015), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1042), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n743), .A2(KEYINPUT53), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n975), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1013), .B2(G2078), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n997), .A2(new_n698), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G171), .ZN(new_n1056));
  NOR4_X1   g631(.A1(new_n1018), .A2(new_n1041), .A3(new_n1049), .A4(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n996), .A2(new_n1005), .A3(new_n1006), .A4(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(new_n1018), .A3(new_n1038), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1021), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G305), .A2(G1981), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G288), .A2(G1976), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1034), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1017), .A2(new_n1008), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1059), .A2(KEYINPUT117), .A3(new_n1038), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1066), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n1041), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n991), .A2(G8), .A3(G168), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1018), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1065), .B1(new_n1073), .B2(KEYINPUT63), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1071), .A2(KEYINPUT63), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1076));
  INV_X1    g651(.A(new_n969), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT123), .B(G2078), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1079), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1053), .A2(G301), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1080), .A2(G301), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT54), .B1(new_n1055), .B2(G171), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1079), .A2(new_n1053), .A3(G301), .A4(new_n1054), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1083), .A2(KEYINPUT54), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n981), .A2(new_n970), .A3(new_n974), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1089), .A2(KEYINPUT122), .B1(new_n1013), .B2(G1996), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1089), .A2(KEYINPUT122), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n558), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n558), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT56), .B(G2072), .Z(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1076), .A2(new_n1097), .A3(new_n979), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n1013), .B2(new_n1098), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n580), .A2(new_n573), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT120), .Z(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n569), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n569), .A2(new_n1105), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT57), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1104), .A2(new_n1108), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1046), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1046), .B2(new_n1111), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1102), .B(new_n1109), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT61), .ZN(new_n1116));
  INV_X1    g691(.A(G1348), .ZN(new_n1117));
  INV_X1    g692(.A(G2067), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n997), .A2(new_n1117), .B1(new_n1019), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n615), .B1(new_n1119), .B2(KEYINPUT60), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1120), .A2(new_n1121), .B1(KEYINPUT60), .B2(new_n1119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1046), .A2(new_n1111), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1112), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1109), .A4(new_n1102), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1096), .A2(new_n1116), .A3(new_n1122), .A4(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1109), .B1(new_n1125), .B2(new_n1102), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1119), .A2(new_n615), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1115), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1086), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1075), .B1(new_n1132), .B2(new_n1003), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1018), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1058), .B(new_n1074), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1012), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n979), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(G1996), .A3(new_n711), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT110), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n734), .A2(G2067), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n729), .A2(new_n1118), .A3(new_n733), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1140), .B(new_n1141), .C1(G1996), .C2(new_n711), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1139), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n816), .A2(new_n819), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n816), .A2(new_n819), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1137), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G290), .B(G1986), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1135), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT127), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1137), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1152), .A2(G1986), .A3(G290), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT48), .Z(new_n1154));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1152), .B1(new_n1157), .B2(new_n1141), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1151), .A2(new_n1156), .B1(new_n1158), .B2(KEYINPUT125), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1158), .A2(KEYINPUT125), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1152), .A2(G1996), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT46), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1137), .B1(new_n1163), .B2(new_n711), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT126), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT47), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1159), .A2(new_n1160), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1150), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g744(.A(new_n865), .ZN(new_n1171));
  NOR2_X1   g745(.A1(new_n959), .A2(new_n960), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n463), .A2(G227), .ZN(new_n1173));
  NAND4_X1  g747(.A1(new_n691), .A2(new_n661), .A3(new_n692), .A4(new_n1173), .ZN(new_n1174));
  NOR3_X1   g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(G308));
  INV_X1    g749(.A(G308), .ZN(G225));
endmodule


