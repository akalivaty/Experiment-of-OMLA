//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n536, new_n537,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n594, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  NOR2_X1   g044(.A1(new_n460), .A2(new_n462), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G124), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT68), .ZN(new_n472));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n461), .B2(G136), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G162));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n478));
  OAI211_X1 g053(.A(G138), .B(new_n462), .C1(new_n458), .C2(new_n459), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n480), .B2(new_n479), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n462), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OR3_X1    g061(.A1(new_n484), .A2(new_n485), .A3(new_n483), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n486), .A2(new_n487), .B1(new_n470), .B2(G126), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n479), .A2(new_n480), .A3(new_n478), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n482), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  INV_X1    g066(.A(G62), .ZN(new_n492));
  OR2_X1    g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G75), .A2(G543), .ZN(new_n496));
  OAI21_X1  g071(.A(G651), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G543), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(new_n499), .A3(G88), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(G50), .A3(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(G303));
  INV_X1    g077(.A(G303), .ZN(G166));
  NAND3_X1  g078(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT7), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n499), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G51), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n499), .A2(G89), .ZN(new_n512));
  NAND2_X1  g087(.A1(G63), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n508), .A2(new_n514), .ZN(G168));
  AOI22_X1  g090(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G52), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n510), .A2(new_n509), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G90), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n506), .A2(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G171));
  AOI22_X1  g100(.A1(new_n498), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n517), .ZN(new_n527));
  INV_X1    g102(.A(new_n522), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n520), .A2(new_n521), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(G81), .B1(new_n531), .B2(G43), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(G153));
  NAND4_X1  g109(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g110(.A1(G1), .A2(G3), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT8), .ZN(new_n537));
  NAND4_X1  g112(.A1(G319), .A2(G483), .A3(G661), .A4(new_n537), .ZN(G188));
  NAND2_X1  g113(.A1(new_n528), .A2(G91), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT9), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n531), .B2(G53), .ZN(new_n541));
  INV_X1    g116(.A(G53), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n506), .A2(KEYINPUT9), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G65), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n511), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  OAI21_X1  g122(.A(G651), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  OAI221_X1 g124(.A(new_n539), .B1(new_n541), .B2(new_n543), .C1(new_n548), .C2(new_n549), .ZN(G299));
  INV_X1    g125(.A(G171), .ZN(G301));
  XNOR2_X1  g126(.A(G168), .B(KEYINPUT72), .ZN(G286));
  OAI211_X1 g127(.A(G49), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n553));
  NOR3_X1   g128(.A1(new_n509), .A2(new_n510), .A3(G74), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(new_n517), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n498), .A2(new_n499), .A3(G87), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT73), .ZN(G288));
  INV_X1    g133(.A(G48), .ZN(new_n559));
  INV_X1    g134(.A(G86), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n506), .A2(new_n559), .B1(new_n522), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  OAI21_X1  g137(.A(G61), .B1(new_n509), .B2(new_n510), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT74), .B1(new_n565), .B2(G651), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  AOI211_X1 g142(.A(new_n567), .B(new_n517), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n562), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n564), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n498), .B2(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n567), .B1(new_n571), .B2(new_n517), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n565), .A2(KEYINPUT74), .A3(G651), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(KEYINPUT75), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n561), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n528), .A2(G85), .B1(new_n531), .B2(G47), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n517), .B2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n528), .A2(G92), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n511), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n531), .B2(G54), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n580), .B1(new_n589), .B2(G868), .ZN(G321));
  XNOR2_X1  g165(.A(G321), .B(KEYINPUT76), .ZN(G284));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G286), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g168(.A(G299), .B(KEYINPUT77), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n592), .ZN(G297));
  XNOR2_X1  g170(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n589), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n533), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g177(.A1(new_n458), .A2(new_n459), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n463), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2100), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n461), .A2(G135), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n470), .A2(G123), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n462), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT79), .B(G2096), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n614), .ZN(G156));
  XOR2_X1   g190(.A(KEYINPUT15), .B(G2435), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2438), .ZN(new_n617));
  XOR2_X1   g192(.A(G2427), .B(G2430), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT82), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n617), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(KEYINPUT14), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G1341), .B(G1348), .Z(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n622), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(G14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT83), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G401));
  INV_X1    g210(.A(KEYINPUT18), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G227));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT84), .Z(new_n655));
  OR2_X1    g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT20), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n653), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n650), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G6), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n575), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT32), .B(G1981), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n674), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n676), .B(new_n672), .C1(new_n575), .C2(new_n671), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n497), .A2(G16), .A3(new_n500), .A4(new_n501), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n679));
  NOR2_X1   g254(.A1(G16), .A2(G22), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AND3_X1   g256(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n679), .B1(new_n678), .B2(new_n681), .ZN(new_n683));
  OAI21_X1  g258(.A(G1971), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT87), .ZN(new_n686));
  INV_X1    g261(.A(G1971), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(KEYINPUT86), .B1(new_n555), .B2(new_n556), .ZN(new_n691));
  OAI21_X1  g266(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n498), .A2(new_n499), .A3(G87), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .A4(new_n553), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(G16), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT33), .B(G1976), .Z(new_n697));
  OR2_X1    g272(.A1(G16), .A2(G23), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n675), .A2(new_n677), .A3(new_n690), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n690), .A2(new_n701), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n677), .A4(new_n675), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n671), .A2(G24), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G290), .B2(G16), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G1986), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n461), .A2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n470), .A2(G119), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n462), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n712), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G25), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n720), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n717), .B(new_n722), .C1(new_n718), .C2(G29), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n710), .A2(new_n711), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n704), .B1(new_n707), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n704), .B(new_n724), .C1(new_n702), .C2(KEYINPUT34), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n703), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT89), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(new_n703), .C1(new_n725), .C2(new_n727), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT36), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT25), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  INV_X1    g314(.A(G127), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n460), .B2(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n741), .A2(G2105), .B1(new_n461), .B2(G139), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT96), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n735), .B1(new_n744), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(G2072), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT98), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n734), .A2(G35), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT100), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n734), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2090), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n671), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n533), .B2(new_n671), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1341), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n461), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n470), .A2(G128), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n462), .A2(G116), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n734), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n671), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT23), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G171), .A2(new_n671), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G5), .B2(new_n671), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n780), .B1(new_n734), .B2(new_n612), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G160), .A2(G29), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G34), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n734), .B1(new_n786), .B2(G34), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n734), .A2(G32), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n470), .A2(G129), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT26), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n463), .A2(G105), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n603), .A2(new_n462), .ZN(new_n797));
  INV_X1    g372(.A(G141), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n791), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT27), .B(G1996), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n789), .A2(new_n790), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n769), .A2(new_n774), .A3(new_n784), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n748), .A2(new_n753), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n802), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  INV_X1    g382(.A(G2078), .ZN(new_n808));
  NAND2_X1  g383(.A1(G164), .A2(G29), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G27), .B2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n808), .ZN(new_n812));
  NOR2_X1   g387(.A1(G168), .A2(new_n671), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n671), .B2(G21), .ZN(new_n814));
  INV_X1    g389(.A(G1966), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n783), .A2(new_n782), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n789), .A2(new_n790), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n816), .B(new_n817), .C1(new_n815), .C2(new_n814), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n811), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G4), .A2(G16), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT91), .Z(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n588), .B2(new_n671), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT93), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT92), .B(G1348), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n745), .A2(new_n746), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT97), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n819), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n805), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n733), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(new_n703), .C1(new_n725), .C2(new_n727), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT90), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n831), .B1(new_n728), .B2(KEYINPUT89), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n732), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n830), .A2(new_n835), .ZN(G311));
  OAI21_X1  g411(.A(KEYINPUT101), .B1(new_n830), .B2(new_n835), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n724), .B1(new_n702), .B2(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT88), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n839), .A2(new_n726), .B1(KEYINPUT34), .B2(new_n702), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT36), .B1(new_n840), .B2(new_n731), .ZN(new_n841));
  INV_X1    g416(.A(new_n732), .ZN(new_n842));
  OAI211_X1 g417(.A(KEYINPUT90), .B(new_n832), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n733), .A4(new_n829), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n837), .A2(new_n845), .ZN(G150));
  NAND2_X1  g421(.A1(new_n589), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n528), .A2(G93), .B1(new_n531), .B2(G55), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT102), .B1(new_n850), .B2(new_n517), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n850), .A2(KEYINPUT102), .A3(new_n517), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n533), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n533), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n848), .B(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT103), .B(G860), .Z(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n854), .A2(new_n862), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n716), .B(KEYINPUT107), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n605), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n461), .A2(G142), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT105), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n462), .A2(KEYINPUT106), .A3(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT106), .B1(new_n462), .B2(G118), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n872), .A2(G2104), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n470), .A2(G130), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n869), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n800), .B(new_n761), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n490), .A2(KEYINPUT104), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n482), .A2(new_n488), .A3(new_n882), .A4(new_n489), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n880), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n744), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n879), .B(new_n886), .C1(new_n743), .C2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n743), .B2(new_n885), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n869), .B(new_n877), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(G160), .B(new_n612), .Z(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(G162), .Z(new_n893));
  OAI21_X1  g468(.A(new_n867), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n887), .A2(KEYINPUT108), .A3(new_n895), .A4(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT40), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(G395));
  XNOR2_X1  g476(.A(new_n588), .B(G299), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(KEYINPUT109), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n857), .B(new_n599), .Z(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n903), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n691), .A2(new_n695), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n575), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(G303), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n917), .B(new_n918), .Z(new_n919));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n912), .B(new_n920), .C1(new_n903), .C2(new_n911), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n914), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n914), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G868), .B2(new_n854), .ZN(G295));
  OAI21_X1  g500(.A(new_n924), .B1(G868), .B2(new_n854), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  NAND3_X1  g503(.A1(G286), .A2(new_n928), .A3(G171), .ZN(new_n929));
  INV_X1    g504(.A(G168), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n930), .B2(G171), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT72), .ZN(new_n932));
  XNOR2_X1  g507(.A(G168), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n933), .B2(G301), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n857), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n857), .B1(new_n929), .B2(new_n934), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n909), .A3(new_n908), .ZN(new_n938));
  INV_X1    g513(.A(new_n919), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n935), .A2(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n903), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n905), .B2(new_n907), .ZN(new_n947));
  INV_X1    g522(.A(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n919), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n943), .A3(new_n942), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n946), .B1(new_n927), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT44), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(KEYINPUT43), .B2(new_n950), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n881), .A2(new_n958), .A3(new_n883), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n464), .A2(new_n468), .A3(G40), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT111), .Z(new_n964));
  INV_X1    g539(.A(new_n800), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(new_n962), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n761), .B(new_n767), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n961), .B2(new_n965), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n964), .A2(new_n965), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n716), .A2(new_n722), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n716), .A2(new_n722), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n968), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(G290), .B(G1986), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n968), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n575), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT119), .Z(new_n983));
  NOR3_X1   g558(.A1(new_n566), .A2(new_n568), .A3(new_n561), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT118), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT49), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n490), .A2(new_n962), .A3(new_n958), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT116), .B(G8), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n986), .B2(KEYINPUT49), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G288), .A2(G1976), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n983), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n988), .B(new_n990), .C1(new_n997), .C2(new_n915), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(KEYINPUT52), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n996), .A3(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(new_n998), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1000), .A2(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n993), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n490), .A2(new_n958), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n490), .A2(new_n1008), .A3(new_n958), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n962), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2090), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n967), .B1(new_n1006), .B2(new_n960), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n958), .A4(new_n883), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1971), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G303), .A2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT113), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  NAND4_X1  g595(.A1(G303), .A2(new_n1020), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1022), .A2(new_n1023), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(KEYINPUT114), .A3(new_n1021), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT115), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1016), .A2(G8), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n995), .A2(new_n991), .B1(new_n1005), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g608(.A(KEYINPUT120), .B1(new_n1005), .B2(new_n1030), .C1(new_n995), .C2(new_n991), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1010), .A2(G2084), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1966), .B1(new_n1012), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G168), .A2(new_n989), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1036), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n930), .B(new_n990), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n990), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1041), .A2(KEYINPUT51), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1043), .A2(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1012), .A2(new_n1013), .A3(new_n808), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1055));
  AOI22_X1  g630(.A1(new_n1054), .A2(new_n1055), .B1(new_n783), .B2(new_n1010), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1012), .A2(new_n1038), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1029), .A2(new_n1026), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n993), .B(new_n1004), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1016), .A2(new_n990), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1051), .A2(new_n1053), .A3(new_n1059), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1001), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(new_n999), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n987), .B2(new_n992), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1060), .B1(new_n989), .B2(new_n1015), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1046), .A2(G286), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1030), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1046), .A2(new_n1073), .A3(G286), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1069), .A2(new_n1030), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1035), .A2(new_n1065), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n966), .A2(new_n962), .A3(new_n1013), .A4(new_n1057), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1056), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1083), .B2(new_n1059), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(G171), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1056), .A2(G301), .A3(new_n1058), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(KEYINPUT54), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1064), .A2(new_n1084), .A3(new_n1087), .A4(new_n1052), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  INV_X1    g664(.A(new_n988), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1010), .A2(new_n1089), .B1(new_n767), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1092), .A2(KEYINPUT122), .A3(new_n588), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n588), .B1(new_n1092), .B2(KEYINPUT122), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(KEYINPUT122), .B2(new_n1092), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1010), .A2(new_n773), .ZN(new_n1098));
  XOR2_X1   g673(.A(G299), .B(KEYINPUT57), .Z(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1012), .A2(new_n1013), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1099), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1012), .A2(new_n1013), .A3(new_n961), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1090), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n533), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1109), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1102), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1097), .A2(new_n1110), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1107), .B1(new_n588), .B2(new_n1091), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1104), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1088), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n980), .B1(new_n1079), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n967), .B(new_n966), .C1(new_n965), .C2(new_n969), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1124), .A2(KEYINPUT126), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(KEYINPUT126), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n963), .B(KEYINPUT111), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT46), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1125), .A2(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT47), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(KEYINPUT125), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(KEYINPUT125), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1129), .B(new_n1130), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1131), .B(KEYINPUT125), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1130), .B1(new_n1136), .B2(new_n1129), .ZN(new_n1137));
  INV_X1    g712(.A(new_n968), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1138), .A2(G1986), .A3(G290), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT48), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1135), .A2(new_n1137), .B1(new_n978), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n761), .A2(G2067), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1123), .A2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g721(.A1(new_n647), .A2(G319), .ZN(new_n1148));
  XOR2_X1   g722(.A(new_n1148), .B(KEYINPUT127), .Z(new_n1149));
  NAND3_X1  g723(.A1(new_n669), .A2(new_n634), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g724(.A(new_n1150), .B1(new_n897), .B2(new_n898), .ZN(new_n1151));
  AND2_X1   g725(.A1(new_n1151), .A2(new_n954), .ZN(G308));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n954), .ZN(G225));
endmodule


