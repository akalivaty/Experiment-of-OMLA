//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OAI211_X1 g003(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n189), .C2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT65), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n188), .B1(new_n191), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n189), .A2(G146), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n198), .A2(new_n193), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n196), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n193), .A2(new_n199), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT0), .B(G128), .Z(new_n205));
  OAI211_X1 g019(.A(new_n204), .B(G125), .C1(new_n205), .C2(new_n187), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G953), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G224), .ZN(new_n209));
  XOR2_X1   g023(.A(new_n207), .B(new_n209), .Z(new_n210));
  XNOR2_X1  g024(.A(G110), .B(G122), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n223), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n218), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(G107), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n229), .A2(new_n232), .A3(new_n236), .A4(new_n233), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(new_n239), .A3(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n227), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n216), .B2(new_n217), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n228), .A2(G107), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n231), .A2(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(G101), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n237), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n224), .A2(KEYINPUT5), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n212), .A3(G116), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n250), .A2(new_n251), .A3(G113), .A4(new_n253), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT5), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(G113), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT84), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n245), .A2(new_n249), .A3(new_n254), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n241), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n211), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n241), .A2(KEYINPUT85), .A3(new_n258), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n241), .A2(new_n211), .A3(new_n258), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n261), .A2(new_n262), .B1(KEYINPUT6), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n210), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G902), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n211), .B(KEYINPUT8), .Z(new_n268));
  NAND3_X1  g082(.A1(new_n250), .A2(G113), .A3(new_n253), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n245), .A2(new_n249), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n245), .A2(new_n254), .A3(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n237), .A2(new_n248), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n270), .B1(new_n273), .B2(KEYINPUT86), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n271), .A2(new_n275), .A3(new_n272), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n268), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n207), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n206), .A2(new_n278), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n281), .A2(new_n282), .A3(new_n202), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n281), .B2(new_n202), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n264), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n267), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT90), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT88), .B(new_n267), .C1(new_n277), .C2(new_n285), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n266), .A2(new_n288), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n290), .B(KEYINPUT91), .Z(new_n295));
  NAND3_X1  g109(.A1(new_n266), .A2(new_n288), .A3(new_n292), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n266), .A2(new_n288), .A3(KEYINPUT89), .A4(new_n292), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G237), .ZN(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT69), .ZN(new_n305));
  OAI211_X1 g119(.A(G214), .B(new_n208), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n189), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(KEYINPUT69), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(G237), .ZN(new_n309));
  AOI21_X1  g123(.A(G953), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(G143), .A3(G214), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT18), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n307), .A2(new_n311), .A3(new_n313), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n196), .A2(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n326), .A3(new_n192), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(G146), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n312), .A2(KEYINPUT92), .A3(new_n314), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n317), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n306), .A2(new_n189), .ZN(new_n333));
  AOI21_X1  g147(.A(G143), .B1(new_n310), .B2(G214), .ZN(new_n334));
  OAI21_X1  g148(.A(G131), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT17), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n307), .A2(new_n337), .A3(new_n311), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n319), .A3(G125), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n322), .B2(new_n340), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(G146), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n312), .A2(KEYINPUT17), .A3(G131), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n228), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n332), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT19), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n323), .A2(new_n326), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n192), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n342), .A2(new_n192), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n335), .A2(new_n338), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n347), .B1(new_n332), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n301), .B1(new_n348), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G475), .A2(G902), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n332), .A2(new_n345), .A3(new_n347), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n331), .A2(new_n318), .A3(new_n329), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n362), .A2(new_n317), .B1(new_n356), .B2(new_n355), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT93), .B(new_n361), .C1(new_n363), .C2(new_n347), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT20), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n348), .A2(new_n358), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G475), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n347), .B1(new_n332), .B2(new_n345), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n348), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n375), .B2(new_n267), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G478), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT15), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT9), .B(G234), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(G217), .A3(new_n208), .ZN(new_n382));
  INV_X1    g196(.A(G134), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n197), .A2(G143), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G128), .B(G143), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT94), .A2(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT94), .A2(G122), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n214), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n214), .A2(G122), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n231), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n391), .A2(G107), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n388), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n231), .A3(new_n393), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n387), .B(new_n383), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(KEYINPUT14), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n214), .A3(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G107), .B1(new_n404), .B2(new_n391), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n399), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n397), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n398), .B1(new_n397), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n382), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT95), .ZN(new_n411));
  INV_X1    g225(.A(new_n382), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n397), .A2(new_n398), .A3(new_n406), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n414), .A3(new_n267), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT96), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n379), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n414), .A3(KEYINPUT96), .A4(new_n267), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(new_n379), .ZN(new_n421));
  INV_X1    g235(.A(G952), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n422), .A2(KEYINPUT97), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(KEYINPUT97), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n208), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(G234), .B2(G237), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  AOI211_X1 g241(.A(new_n267), .B(new_n208), .C1(G234), .C2(G237), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n372), .A2(new_n377), .A3(new_n421), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G214), .B1(G237), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n300), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT11), .B1(new_n383), .B2(G137), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT11), .ZN(new_n437));
  INV_X1    g251(.A(G137), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(G134), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT64), .B1(new_n438), .B2(G134), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT64), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n383), .A3(G137), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n440), .A2(G131), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n441), .A2(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n436), .A2(new_n439), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n337), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n435), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n204), .B1(new_n205), .B2(new_n187), .ZN(new_n450));
  OAI21_X1  g264(.A(G131), .B1(new_n440), .B2(new_n444), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n337), .A3(new_n447), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT67), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n383), .A2(G137), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n438), .A2(G134), .ZN(new_n456));
  OAI21_X1  g270(.A(G131), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT1), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(G143), .B2(new_n192), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n197), .B1(new_n459), .B2(KEYINPUT65), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n187), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n452), .B(new_n457), .C1(new_n464), .C2(new_n200), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n465), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n243), .A2(new_n244), .B1(new_n216), .B2(new_n217), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n310), .A2(G210), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT27), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(G101), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n452), .A2(new_n457), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n463), .A2(G128), .A3(new_n190), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n200), .B1(new_n479), .B2(new_n188), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n450), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n451), .B2(new_n452), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n227), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT68), .B1(new_n478), .B2(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n195), .A2(new_n201), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n452), .A4(new_n457), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n454), .A2(new_n470), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n450), .B1(new_n445), .B2(new_n448), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n465), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT72), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n227), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n473), .A2(new_n477), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n454), .A2(KEYINPUT30), .A3(new_n486), .A4(new_n489), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n470), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n490), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT74), .ZN(new_n505));
  INV_X1    g319(.A(new_n477), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n454), .A2(new_n486), .A3(new_n489), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n509), .A2(new_n470), .B1(new_n500), .B2(new_n502), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT74), .B1(new_n510), .B2(new_n477), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n498), .A2(new_n499), .A3(new_n507), .A4(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n227), .B1(new_n466), .B2(new_n467), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n513), .B2(new_n469), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n227), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n472), .B1(new_n515), .B2(new_n490), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n506), .A2(new_n499), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G472), .ZN(new_n521));
  INV_X1    g335(.A(new_n496), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n493), .B1(new_n492), .B2(new_n227), .ZN(new_n523));
  AOI211_X1 g337(.A(KEYINPUT72), .B(new_n470), .C1(new_n465), .C2(new_n491), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n522), .B1(new_n525), .B2(new_n490), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n506), .B1(new_n526), .B2(new_n514), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n500), .A2(new_n502), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n490), .A2(new_n477), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT31), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT70), .ZN(new_n531));
  OR3_X1    g345(.A1(new_n528), .A2(KEYINPUT31), .A3(new_n529), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n503), .A2(new_n477), .A3(new_n490), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT31), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n527), .A2(new_n531), .A3(new_n532), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT32), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n521), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n212), .B2(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n212), .A2(G128), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(G110), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n197), .A2(G119), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G110), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT75), .B1(new_n546), .B2(G110), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT76), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n549), .A2(new_n555), .A3(new_n558), .A4(new_n553), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n354), .A2(new_n327), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n343), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n551), .A2(new_n552), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G110), .B2(new_n546), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT22), .B(G137), .ZN(new_n568));
  INV_X1    g382(.A(G221), .ZN(new_n569));
  INV_X1    g383(.A(G234), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n569), .A2(new_n570), .A3(G953), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n568), .B(new_n571), .Z(new_n572));
  NAND3_X1  g386(.A1(new_n563), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n572), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n561), .B1(new_n557), .B2(new_n559), .ZN(new_n575));
  INV_X1    g389(.A(new_n567), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G217), .B1(new_n570), .B2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n267), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT78), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT78), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n573), .A2(new_n577), .A3(new_n583), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n573), .A2(new_n577), .A3(new_n586), .A4(new_n267), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n573), .A2(new_n267), .A3(new_n577), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n578), .B1(new_n588), .B2(KEYINPUT25), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n569), .B1(new_n381), .B2(new_n267), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n267), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT79), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n237), .A2(new_n248), .A3(KEYINPUT10), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n480), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n487), .A2(new_n597), .A3(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n240), .A2(new_n450), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n461), .A2(G128), .B1(new_n193), .B2(new_n199), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n237), .B(new_n248), .C1(new_n602), .C2(new_n200), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n600), .A2(new_n238), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n449), .A2(new_n605), .A3(new_n453), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n449), .B2(new_n453), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n599), .B(new_n604), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n449), .A2(new_n453), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT83), .B(new_n609), .C1(new_n599), .C2(new_n604), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT83), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT79), .B1(new_n487), .B2(new_n597), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n480), .A2(new_n594), .A3(new_n595), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n604), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n609), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n608), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(G110), .B(G140), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n208), .A2(G227), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n195), .A2(new_n272), .A3(new_n201), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n603), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n449), .A3(new_n453), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT12), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n451), .A2(new_n452), .ZN(new_n627));
  NOR2_X1   g441(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n628));
  AND2_X1   g442(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n623), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n620), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n608), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n621), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n593), .B1(new_n635), .B2(new_n592), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n608), .A2(new_n631), .A3(KEYINPUT82), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT82), .B1(new_n608), .B2(new_n631), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n620), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n608), .A2(new_n632), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n234), .A2(G101), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n450), .B(new_n240), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n603), .A2(new_n601), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n596), .B2(new_n598), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT83), .B1(new_n646), .B2(new_n609), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n614), .A2(new_n611), .A3(new_n615), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n639), .A2(G469), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n591), .B1(new_n636), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n434), .A2(new_n541), .A3(new_n590), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G101), .ZN(G3));
  NAND2_X1  g468(.A1(new_n536), .A2(new_n267), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT98), .B1(new_n655), .B2(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n536), .A2(new_n538), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n531), .A2(new_n535), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n533), .A2(KEYINPUT31), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n473), .A2(new_n497), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n506), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G472), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n656), .B1(new_n664), .B2(KEYINPUT98), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n296), .A2(new_n290), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n433), .B1(new_n666), .B2(new_n293), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n430), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n409), .A2(new_n414), .A3(KEYINPUT33), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT33), .B1(new_n409), .B2(new_n414), .ZN(new_n670));
  OAI211_X1 g484(.A(G478), .B(new_n267), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n415), .A2(new_n378), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n370), .B1(new_n365), .B2(KEYINPUT20), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n376), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n632), .B1(new_n649), .B2(new_n608), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n592), .B(new_n267), .C1(new_n677), .C2(new_n633), .ZN(new_n678));
  INV_X1    g492(.A(new_n593), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n651), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n591), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n680), .A2(new_n590), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n665), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT34), .B(G104), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G6));
  XNOR2_X1  g499(.A(new_n365), .B(KEYINPUT20), .ZN(new_n686));
  INV_X1    g500(.A(new_n421), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n377), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n668), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n665), .A2(new_n682), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT99), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT35), .B(G107), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NAND2_X1  g507(.A1(new_n296), .A2(new_n297), .ZN(new_n694));
  INV_X1    g508(.A(new_n295), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n299), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n293), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n420), .A2(new_n379), .ZN(new_n698));
  INV_X1    g512(.A(new_n417), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n430), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n376), .A3(new_n674), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n652), .A2(new_n697), .A3(new_n432), .A4(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n663), .B1(new_n536), .B2(new_n267), .ZN(new_n703));
  INV_X1    g517(.A(new_n538), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n658), .B2(new_n661), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT98), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT98), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n662), .B2(new_n663), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n589), .A2(new_n587), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n575), .A2(KEYINPUT36), .A3(new_n576), .A4(new_n574), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n563), .B2(new_n567), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n580), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n708), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n702), .B1(new_n716), .B2(KEYINPUT100), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n665), .A2(new_n718), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT37), .B(G110), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G12));
  NAND3_X1  g536(.A1(new_n680), .A2(new_n681), .A3(new_n715), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n666), .A2(new_n293), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n432), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(G900), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n426), .B1(new_n727), .B2(new_n428), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n688), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n729), .A3(new_n541), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G128), .ZN(G30));
  XOR2_X1   g545(.A(new_n728), .B(KEYINPUT39), .Z(new_n732));
  AND2_X1   g546(.A1(new_n652), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT40), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n300), .B(KEYINPUT38), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n510), .A2(new_n506), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n515), .A2(new_n506), .A3(new_n490), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n267), .ZN(new_n738));
  OAI21_X1  g552(.A(G472), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n539), .B2(new_n540), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n421), .B1(new_n372), .B2(new_n377), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n709), .A2(new_n714), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n432), .A3(new_n743), .ZN(new_n744));
  OR4_X1    g558(.A1(new_n734), .A2(new_n735), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G143), .ZN(G45));
  INV_X1    g560(.A(new_n728), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n673), .B(new_n747), .C1(new_n674), .C2(new_n376), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n726), .A2(new_n541), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G146), .ZN(G48));
  INV_X1    g565(.A(new_n590), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n657), .A2(KEYINPUT32), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n752), .B1(new_n755), .B2(new_n521), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n592), .A2(KEYINPUT101), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n677), .A2(new_n633), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(G902), .ZN(new_n759));
  INV_X1    g573(.A(new_n757), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n635), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n681), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n756), .A2(new_n676), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(KEYINPUT41), .B(G113), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G15));
  NAND3_X1  g580(.A1(new_n756), .A2(new_n689), .A3(new_n763), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G116), .ZN(G18));
  NOR2_X1   g582(.A1(new_n725), .A2(new_n762), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n541), .A3(new_n701), .A4(new_n715), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G119), .ZN(G21));
  NAND2_X1  g585(.A1(new_n742), .A2(new_n667), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n772), .A2(new_n429), .A3(new_n762), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n532), .A2(new_n530), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n506), .B1(new_n514), .B2(new_n516), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n704), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n752), .A2(new_n703), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NOR3_X1   g593(.A1(new_n703), .A2(new_n743), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n748), .A2(KEYINPUT102), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n372), .A2(new_n377), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT102), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n673), .A4(new_n747), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n769), .A2(new_n780), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G125), .ZN(G27));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n300), .A2(new_n432), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT103), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n651), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n639), .A2(KEYINPUT103), .A3(G469), .A4(new_n650), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n678), .A3(new_n679), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n681), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT104), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(KEYINPUT104), .A3(new_n681), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n756), .A2(new_n789), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n784), .A2(new_n781), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n787), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n796), .A2(new_n797), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n541), .A2(new_n590), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n788), .ZN(new_n803));
  INV_X1    g617(.A(new_n799), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT42), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G131), .ZN(G33));
  XOR2_X1   g621(.A(new_n729), .B(KEYINPUT105), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n803), .A3(new_n801), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G134), .ZN(G36));
  AND2_X1   g624(.A1(new_n639), .A2(new_n650), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT45), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT45), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(G469), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n679), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n816), .B1(new_n592), .B2(new_n635), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n681), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n732), .A3(new_n789), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT106), .ZN(new_n822));
  INV_X1    g636(.A(new_n673), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n782), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT43), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT107), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n665), .A2(new_n743), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n826), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n821), .B1(new_n831), .B2(KEYINPUT44), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT108), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n831), .B2(KEYINPUT44), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT44), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G137), .ZN(G39));
  XOR2_X1   g651(.A(new_n819), .B(KEYINPUT47), .Z(new_n838));
  NOR4_X1   g652(.A1(new_n541), .A2(new_n788), .A3(new_n590), .A4(new_n748), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT109), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(KEYINPUT110), .B(G140), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(G42));
  NAND3_X1  g657(.A1(new_n706), .A2(new_n682), .A3(new_n708), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n433), .B1(new_n696), .B2(new_n293), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n782), .A2(new_n421), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n430), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n717), .B2(new_n719), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n675), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(KEYINPUT112), .B(new_n673), .C1(new_n674), .C2(new_n376), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n845), .A2(new_n430), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  OAI22_X1  g667(.A1(new_n844), .A2(new_n853), .B1(new_n802), .B2(new_n702), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n653), .B(new_n856), .C1(new_n844), .C2(new_n853), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n849), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n849), .A2(new_n855), .A3(new_n857), .A4(KEYINPUT114), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n686), .A2(new_n377), .A3(new_n421), .A4(new_n747), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT115), .ZN(new_n864));
  INV_X1    g678(.A(new_n723), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n541), .A3(new_n865), .A4(new_n789), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n801), .A2(new_n780), .A3(new_n804), .A4(new_n789), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n809), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n726), .B(new_n541), .C1(new_n729), .C2(new_n749), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n709), .A2(new_n714), .A3(new_n747), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n742), .A2(new_n667), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n681), .A3(new_n740), .A4(new_n793), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n873), .A3(new_n785), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n870), .A2(new_n873), .A3(new_n785), .A4(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n764), .A2(new_n767), .A3(new_n770), .A4(new_n778), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n878), .A2(new_n806), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n862), .A2(new_n869), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(new_n806), .A3(KEYINPUT53), .A4(new_n879), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n868), .B1(new_n860), .B2(new_n861), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(KEYINPUT117), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n888), .B(new_n868), .C1(new_n860), .C2(new_n861), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n878), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n881), .A2(new_n882), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n881), .B1(new_n882), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n825), .A2(new_n426), .A3(new_n777), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n759), .A2(new_n761), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n681), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n789), .B(new_n897), .C1(new_n838), .C2(new_n899), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n426), .A2(new_n825), .A3(new_n763), .A4(new_n789), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n780), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n590), .A2(new_n426), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n740), .A2(new_n788), .A3(new_n762), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(new_n377), .A3(new_n372), .A4(new_n823), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n735), .A2(new_n433), .A3(new_n763), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n897), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT50), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n900), .A2(new_n914), .A3(KEYINPUT51), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT51), .B1(new_n900), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n901), .A2(new_n756), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT48), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n897), .A2(new_n769), .ZN(new_n919));
  INV_X1    g733(.A(new_n675), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n425), .B1(new_n904), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n891), .A2(new_n896), .A3(new_n915), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n898), .B(KEYINPUT49), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n590), .A2(new_n681), .A3(new_n432), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n927), .A2(new_n782), .A3(new_n823), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n926), .A2(new_n735), .A3(new_n741), .A4(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT111), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G75));
  NOR2_X1   g745(.A1(new_n208), .A2(G952), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n862), .A2(new_n869), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n888), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n886), .A2(KEYINPUT117), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n935), .A3(new_n885), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n267), .B1(new_n936), .B2(new_n883), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n937), .B2(new_n290), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n263), .A2(new_n265), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n210), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n937), .A2(new_n695), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT56), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n932), .B(new_n942), .C1(new_n943), .C2(new_n947), .ZN(G51));
  OR3_X1    g762(.A1(new_n890), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT120), .B1(new_n890), .B2(KEYINPUT54), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n593), .B(KEYINPUT57), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n758), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n937), .A2(G469), .A3(new_n813), .A4(new_n812), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n932), .B1(new_n956), .B2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n359), .A2(new_n364), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n932), .ZN(G60));
  INV_X1    g777(.A(new_n932), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n891), .B2(new_n896), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n669), .A2(new_n670), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(new_n966), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n952), .B2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n890), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n713), .ZN(new_n977));
  OAI211_X1 g791(.A(KEYINPUT61), .B(new_n964), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n573), .A2(new_n577), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT122), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT122), .ZN(new_n981));
  INV_X1    g795(.A(new_n979), .ZN(new_n982));
  AOI211_X1 g796(.A(new_n981), .B(new_n982), .C1(new_n890), .C2(new_n975), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n978), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n974), .B1(new_n936), .B2(new_n883), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n932), .B1(new_n987), .B2(new_n713), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n890), .B2(new_n975), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT123), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n964), .B1(new_n976), .B2(new_n977), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n985), .B1(new_n994), .B2(new_n989), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n989), .B(KEYINPUT122), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n993), .B(new_n995), .C1(new_n996), .C2(new_n978), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n992), .A2(new_n997), .ZN(G66));
  INV_X1    g812(.A(G224), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n427), .B2(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n862), .A2(new_n879), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n939), .B1(G898), .B2(new_n208), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G69));
  AOI21_X1  g818(.A(new_n208), .B1(G227), .B2(G900), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n802), .A2(new_n772), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n820), .A2(new_n732), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n870), .A2(new_n785), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1008), .A2(new_n809), .A3(new_n1010), .ZN(new_n1011));
  AND4_X1   g825(.A1(new_n806), .A2(new_n836), .A3(new_n841), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n208), .ZN(new_n1013));
  INV_X1    g827(.A(new_n492), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n500), .B1(KEYINPUT30), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT124), .Z(new_n1016));
  NAND2_X1  g830(.A1(new_n350), .A2(new_n351), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1016), .B(new_n1017), .Z(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(G900), .B2(G953), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n745), .A2(new_n1010), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT62), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n838), .B2(new_n840), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n851), .A2(new_n852), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n803), .B(new_n733), .C1(new_n846), .C2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n836), .A2(KEYINPUT126), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(KEYINPUT126), .B1(new_n836), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1024), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1030), .A2(new_n208), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1018), .B(KEYINPUT125), .Z(new_n1032));
  OAI211_X1 g846(.A(new_n1006), .B(new_n1021), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1032), .B1(new_n1030), .B2(new_n208), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1021), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1005), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1033), .A2(new_n1036), .ZN(G72));
  NOR2_X1   g851(.A1(new_n894), .A2(new_n895), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n511), .A2(new_n533), .A3(new_n507), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT127), .Z(new_n1043));
  NOR2_X1   g857(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1041), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1045), .B1(new_n1012), .B2(new_n1001), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n510), .A2(new_n506), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n964), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n862), .A2(new_n879), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1041), .B1(new_n1030), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g864(.A(new_n1044), .B(new_n1048), .C1(new_n736), .C2(new_n1050), .ZN(G57));
endmodule


