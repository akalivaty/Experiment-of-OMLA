//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT72), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n214), .B1(new_n210), .B2(new_n211), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G190gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(KEYINPUT23), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n217), .B2(G190gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(KEYINPUT23), .B2(new_n220), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT25), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n230), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G183gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n237), .A3(new_n228), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT28), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT28), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n228), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n228), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n250), .B1(new_n249), .B2(new_n252), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n244), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n222), .A2(new_n225), .A3(KEYINPUT25), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n231), .B1(new_n230), .B2(new_n221), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n233), .A2(new_n256), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(KEYINPUT29), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n226), .A2(new_n232), .ZN(new_n264));
  NOR3_X1   g063(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n248), .ZN(new_n266));
  INV_X1    g065(.A(new_n245), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT66), .B1(new_n268), .B2(new_n251), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n243), .B1(new_n269), .B2(new_n253), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n263), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n216), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n233), .A2(new_n256), .A3(new_n260), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(new_n261), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n264), .A2(new_n270), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n273), .A2(new_n276), .B1(new_n277), .B2(new_n261), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n272), .B1(new_n278), .B2(new_n216), .ZN(new_n279));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT74), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n273), .A2(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(new_n261), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n216), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n271), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n213), .A2(new_n215), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n287), .A2(new_n290), .A3(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT30), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n287), .A2(new_n290), .A3(new_n298), .A4(new_n283), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n294), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n295), .B1(new_n294), .B2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G127gat), .ZN(new_n306));
  INV_X1    g105(.A(G127gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(KEYINPUT1), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n312), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(G113gat), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT67), .B1(new_n312), .B2(G113gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n306), .A2(new_n308), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g119(.A(new_n318), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n315), .A2(new_n314), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(new_n313), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n311), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT2), .ZN(new_n331));
  XNOR2_X1  g130(.A(G155gat), .B(G162gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n329), .B(new_n331), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n333), .ZN(new_n338));
  XNOR2_X1  g137(.A(G141gat), .B(G148gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(G155gat), .B2(G162gat), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n304), .B1(new_n326), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n334), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n334), .A2(new_n342), .A3(new_n348), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n343), .A2(KEYINPUT3), .B1(new_n323), .B2(new_n311), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n323), .A2(new_n334), .A3(new_n342), .A4(new_n311), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(new_n304), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n344), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n319), .A2(new_n343), .A3(KEYINPUT77), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT77), .B1(new_n319), .B2(new_n343), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n353), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n358), .B(KEYINPUT39), .C1(new_n357), .C2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G1gat), .B(G29gat), .Z(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n362), .B(new_n367), .C1(KEYINPUT39), .C2(new_n358), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n343), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n320), .A2(new_n325), .A3(KEYINPUT4), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n357), .B1(new_n353), .B2(new_n304), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n361), .A2(new_n357), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT5), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n344), .A2(new_n354), .A3(new_n352), .A4(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(new_n367), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n368), .B2(new_n369), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n303), .A2(new_n370), .A3(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n279), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n279), .A2(KEYINPUT86), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT37), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n282), .B1(new_n279), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT38), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n376), .A2(new_n367), .A3(new_n378), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT79), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n376), .A2(new_n404), .A3(new_n367), .A4(new_n378), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n400), .B1(new_n406), .B2(new_n380), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n390), .B1(new_n278), .B2(new_n289), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n288), .A2(new_n216), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT38), .B(new_n283), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n389), .A2(new_n410), .B1(new_n279), .B2(new_n283), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n398), .A3(new_n407), .A4(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n275), .B1(new_n347), .B2(new_n349), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n289), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n212), .A2(new_n274), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n371), .B1(new_n417), .B2(new_n345), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n212), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n345), .B1(new_n420), .B2(KEYINPUT29), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n421), .B2(new_n343), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n415), .B2(new_n289), .ZN(new_n423));
  INV_X1    g222(.A(G22gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n419), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n419), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n413), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n419), .A2(new_n423), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G22gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n419), .A2(new_n423), .A3(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(KEYINPUT82), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT31), .B(G50gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n427), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n413), .B(new_n434), .C1(new_n425), .C2(new_n426), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n382), .A2(new_n412), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n273), .A2(new_n320), .A3(new_n325), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n326), .A2(new_n233), .A3(new_n256), .A4(new_n260), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(G227gat), .A3(G233gat), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(KEYINPUT32), .ZN(new_n446));
  XOR2_X1   g245(.A(G15gat), .B(G43gat), .Z(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT69), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT70), .ZN(new_n449));
  XOR2_X1   g248(.A(G71gat), .B(G99gat), .Z(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT32), .B(new_n443), .C1(new_n453), .C2(new_n444), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n442), .ZN(new_n457));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n459), .B2(KEYINPUT71), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n461), .B(KEYINPUT34), .C1(new_n457), .C2(new_n458), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n452), .B(new_n454), .C1(new_n460), .C2(new_n462), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n403), .A2(new_n405), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n399), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n379), .A2(new_n367), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n284), .A2(new_n293), .B1(new_n297), .B2(new_n299), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n400), .A4(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n476), .B(new_n400), .C1(new_n406), .C2(new_n380), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n438), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n440), .A2(new_n470), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT88), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n303), .B2(new_n407), .ZN(new_n484));
  INV_X1    g283(.A(new_n302), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n295), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n407), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT88), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n464), .A2(new_n436), .A3(new_n465), .A4(new_n437), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AND4_X1   g291(.A1(new_n464), .A2(new_n436), .A3(new_n465), .A4(new_n437), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n479), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n482), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT104), .ZN(new_n498));
  XOR2_X1   g297(.A(G134gat), .B(G162gat), .Z(new_n499));
  XOR2_X1   g298(.A(G43gat), .B(G50gat), .Z(new_n500));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  INV_X1    g304(.A(G36gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n507), .A2(new_n508), .B1(G29gat), .B2(G36gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n502), .A2(new_n503), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n509), .A2(new_n511), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n502), .A2(new_n509), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n519), .A3(new_n516), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT99), .B(G92gat), .Z(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(G85gat), .ZN(new_n523));
  XOR2_X1   g322(.A(G99gat), .B(G106gat), .Z(new_n524));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n524), .A2(new_n525), .B1(KEYINPUT8), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(KEYINPUT98), .A3(KEYINPUT7), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n531), .B(new_n532), .C1(KEYINPUT7), .C2(new_n528), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n523), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n524), .A2(new_n525), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n537), .A2(new_n523), .A3(new_n527), .A4(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n539), .ZN(new_n542));
  AND2_X1   g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT41), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n539), .B1(new_n518), .B2(new_n520), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n547), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n543), .A2(KEYINPUT41), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n549), .B2(new_n551), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n499), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n549), .A2(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n552), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n559));
  INV_X1    g358(.A(new_n499), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563));
  XNOR2_X1  g362(.A(G127gat), .B(G155gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n570), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT96), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT97), .Z(new_n581));
  AND3_X1   g380(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n577), .B2(new_n579), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n565), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n579), .ZN(new_n585));
  INV_X1    g384(.A(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n588), .A3(new_n564), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n584), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n584), .B2(new_n589), .ZN(new_n593));
  INV_X1    g392(.A(G1gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G15gat), .B(G22gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n596), .B2(KEYINPUT92), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT16), .B1(new_n594), .B2(KEYINPUT92), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G8gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n574), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(KEYINPUT21), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n592), .A2(new_n593), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n582), .A2(new_n583), .A3(new_n565), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n564), .B1(new_n587), .B2(new_n588), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n590), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n584), .A2(new_n589), .A3(new_n591), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n563), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n603), .B1(new_n592), .B2(new_n593), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n605), .A3(new_n609), .ZN(new_n613));
  INV_X1    g412(.A(new_n563), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n562), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT102), .ZN(new_n618));
  XOR2_X1   g417(.A(G176gat), .B(G204gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n539), .A2(new_n602), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n536), .A2(new_n574), .A3(new_n538), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT101), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627));
  AOI211_X1 g426(.A(new_n627), .B(new_n624), .C1(new_n621), .C2(new_n622), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n630), .A3(new_n622), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n625), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n620), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  INV_X1    g434(.A(new_n620), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n635), .B(new_n636), .C1(new_n626), .C2(new_n628), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n637), .A3(KEYINPUT103), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT103), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n498), .B1(new_n616), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT90), .ZN(new_n644));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G8gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n600), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n521), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n601), .A2(new_n517), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n653), .A2(KEYINPUT18), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n654), .B(KEYINPUT13), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n516), .A3(new_n514), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n655), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT93), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI211_X1 g461(.A(KEYINPUT93), .B(new_n658), .C1(new_n659), .C2(new_n655), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n656), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n601), .B1(new_n518), .B2(new_n520), .ZN(new_n665));
  INV_X1    g464(.A(new_n655), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT18), .B1(new_n667), .B2(new_n654), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n650), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n654), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n660), .B(new_n661), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n656), .A4(new_n649), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n614), .B1(new_n612), .B2(new_n613), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n639), .A2(new_n640), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n678), .A2(KEYINPUT104), .A3(new_n562), .A4(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n642), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n497), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n488), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n594), .ZN(G1324gat));
  NOR2_X1   g483(.A1(new_n682), .A2(new_n487), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT42), .B1(new_n685), .B2(new_n651), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g487(.A(KEYINPUT42), .B(new_n686), .S(new_n688), .Z(G1325gat));
  INV_X1    g488(.A(new_n466), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n682), .A2(G15gat), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n682), .B2(new_n470), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1326gat));
  NAND3_X1  g492(.A1(new_n497), .A2(new_n438), .A3(new_n681), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT105), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  AOI21_X1  g496(.A(new_n562), .B1(new_n482), .B2(new_n496), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n556), .A2(new_n561), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n492), .A2(new_n495), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n482), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n492), .B2(new_n495), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n699), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n669), .A2(new_n674), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n678), .A2(new_n641), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n488), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n698), .A2(new_n709), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n505), .A3(new_n407), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(G1328gat));
  NOR2_X1   g515(.A1(new_n487), .A2(G36gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n710), .B2(new_n487), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  INV_X1    g527(.A(new_n470), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n707), .A2(new_n728), .A3(new_n729), .A4(new_n709), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n706), .A2(new_n700), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n731), .A2(new_n729), .A3(new_n709), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n727), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n698), .A2(new_n727), .A3(new_n466), .A4(new_n709), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT109), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n733), .B2(G43gat), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n735), .A2(new_n739), .B1(new_n740), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g540(.A1(new_n731), .A2(new_n438), .A3(new_n709), .A4(new_n732), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G50gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n439), .A2(G50gat), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT111), .Z(new_n745));
  NAND2_X1  g544(.A1(new_n712), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n496), .A2(KEYINPUT107), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n482), .A3(new_n703), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n616), .A2(new_n675), .A3(new_n679), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n407), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g554(.A(new_n487), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT112), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n757), .B(new_n759), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n753), .A2(new_n761), .A3(new_n466), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n753), .A2(new_n729), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(new_n761), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n753), .A2(new_n438), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g568(.A1(new_n678), .A2(new_n675), .A3(new_n679), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n707), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n407), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G85gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n678), .A2(new_n675), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n701), .B(new_n774), .C1(new_n704), .C2(new_n705), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n751), .A2(KEYINPUT51), .A3(new_n701), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n679), .A2(new_n488), .A3(G85gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n731), .A2(new_n303), .A3(new_n732), .A4(new_n770), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n522), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n487), .A2(new_n679), .A3(G92gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n784), .B(new_n785), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  AND4_X1   g589(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT52), .A4(new_n789), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(G1337gat));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n779), .A2(new_n793), .A3(new_n466), .A4(new_n641), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n771), .A2(new_n729), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(G1338gat));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n679), .A2(new_n439), .A3(G106gat), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n780), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n731), .A2(new_n438), .A3(new_n732), .A4(new_n770), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n798), .B(KEYINPUT114), .Z(new_n803));
  AOI22_X1  g602(.A1(G106gat), .A2(new_n801), .B1(new_n779), .B2(new_n803), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n800), .A2(new_n802), .B1(new_n804), .B2(new_n797), .ZN(G1339gat));
  NAND4_X1  g604(.A1(new_n678), .A2(new_n708), .A3(new_n562), .A4(new_n679), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n616), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(KEYINPUT115), .A3(new_n708), .A4(new_n679), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n678), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n631), .A2(new_n632), .A3(new_n625), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT54), .B(new_n635), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n636), .B1(new_n633), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n821), .A2(new_n675), .A3(new_n637), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n659), .A2(new_n655), .A3(new_n658), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n667), .B2(new_n654), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n825), .A2(KEYINPUT117), .A3(new_n648), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n825), .B2(new_n648), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n674), .C1(new_n639), .C2(new_n640), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n701), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n821), .A2(new_n637), .A3(new_n822), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n701), .A3(new_n674), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n812), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n488), .B1(new_n811), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n493), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n487), .A3(new_n675), .ZN(new_n840));
  INV_X1    g639(.A(G113gat), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n835), .A2(new_n487), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n493), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n708), .A2(new_n841), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n840), .A2(new_n841), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n487), .A3(new_n641), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n679), .A2(new_n312), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n846), .A2(new_n312), .B1(new_n843), .B2(new_n847), .ZN(G1341gat));
  NAND2_X1  g647(.A1(new_n839), .A2(new_n487), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n678), .A2(new_n307), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n843), .A2(new_n678), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n849), .A2(new_n850), .B1(new_n307), .B2(new_n851), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n303), .A2(new_n562), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G134gat), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n303), .A2(new_n562), .A3(G134gat), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n839), .B2(new_n856), .ZN(new_n857));
  AND4_X1   g656(.A1(KEYINPUT56), .A2(new_n837), .A3(new_n838), .A4(new_n856), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(G1343gat));
  NAND3_X1  g658(.A1(new_n470), .A2(new_n407), .A3(new_n487), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n811), .A2(new_n834), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n438), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n438), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(G141gat), .A3(new_n675), .ZN(new_n867));
  INV_X1    g666(.A(G141gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n470), .A2(new_n438), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n842), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n871), .B2(new_n708), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n873), .B(new_n874), .ZN(G1344gat));
  XOR2_X1   g674(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n876));
  INV_X1    g675(.A(new_n860), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n863), .B(new_n439), .C1(new_n811), .C2(new_n834), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n642), .A2(new_n680), .A3(new_n708), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n834), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n438), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n641), .B(new_n877), .C1(new_n878), .C2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G148gat), .B1(new_n882), .B2(KEYINPUT120), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n822), .A2(new_n637), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n708), .A3(new_n820), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n674), .B1(new_n826), .B2(new_n827), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n679), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n562), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n833), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n678), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n642), .A2(new_n708), .A3(new_n680), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n438), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n863), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n679), .B1(new_n894), .B2(new_n865), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n884), .B1(new_n895), .B2(new_n877), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n876), .B1(new_n883), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(G148gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .ZN(new_n899));
  INV_X1    g698(.A(new_n866), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n679), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n842), .A2(new_n898), .A3(new_n641), .A4(new_n870), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1345gat));
  INV_X1    g703(.A(G155gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n866), .B2(new_n678), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n871), .A2(G155gat), .A3(new_n812), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT121), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT121), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1346gat));
  INV_X1    g709(.A(G162gat), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n866), .A2(new_n701), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(KEYINPUT122), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(KEYINPUT122), .B2(new_n912), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n835), .A2(new_n911), .A3(new_n853), .A4(new_n870), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  AOI21_X1  g715(.A(new_n407), .B1(new_n811), .B2(new_n834), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(new_n493), .A3(new_n303), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n708), .A2(G169gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n487), .A2(new_n407), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT124), .A3(new_n466), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT124), .B1(new_n923), .B2(new_n466), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(new_n438), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n861), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n675), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G169gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n921), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n921), .A2(new_n932), .A3(new_n922), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1348gat));
  INV_X1    g733(.A(G176gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n935), .A3(new_n641), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n927), .A2(new_n641), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n935), .ZN(G1349gat));
  AOI21_X1  g737(.A(new_n234), .B1(new_n927), .B2(new_n678), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n678), .A2(new_n240), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n918), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g741(.A1(new_n918), .A2(new_n228), .A3(new_n701), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n701), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(G190gat), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT61), .B(new_n228), .C1(new_n927), .C2(new_n701), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n948), .B(new_n949), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n869), .A2(new_n487), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n917), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n675), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n470), .A2(new_n923), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n894), .B2(new_n865), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n675), .A2(G197gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  NOR3_X1   g758(.A1(new_n953), .A2(G204gat), .A3(new_n679), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n895), .A2(new_n470), .A3(new_n923), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G204gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n954), .A2(new_n204), .A3(new_n678), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n957), .A2(new_n678), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n966), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n205), .A3(new_n701), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n957), .A2(new_n701), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n972), .B2(new_n205), .ZN(G1355gat));
endmodule


