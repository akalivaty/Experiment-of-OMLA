

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813;

  BUF_X1 U377 ( .A(n737), .Z(n356) );
  AND2_X1 U378 ( .A1(n672), .A2(n671), .ZN(n425) );
  INV_X1 U379 ( .A(G953), .ZN(n805) );
  AND2_X2 U380 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X2 U381 ( .A(n380), .B(n379), .ZN(n653) );
  NOR2_X2 U382 ( .A1(n644), .A2(n760), .ZN(n380) );
  XNOR2_X2 U383 ( .A(n633), .B(n632), .ZN(n705) );
  NOR2_X2 U384 ( .A1(n676), .A2(n675), .ZN(n428) );
  XNOR2_X2 U385 ( .A(n500), .B(KEYINPUT69), .ZN(n547) );
  NOR2_X1 U386 ( .A1(n801), .A2(n473), .ZN(n478) );
  AND2_X1 U387 ( .A1(n459), .A2(n365), .ZN(n458) );
  AND2_X1 U388 ( .A1(n463), .A2(n590), .ZN(n572) );
  AND2_X1 U389 ( .A1(n441), .A2(n439), .ZN(n438) );
  XNOR2_X1 U390 ( .A(n391), .B(KEYINPUT41), .ZN(n779) );
  AND2_X1 U391 ( .A1(n625), .A2(n627), .ZN(n444) );
  XNOR2_X1 U392 ( .A(n427), .B(KEYINPUT112), .ZN(n593) );
  OR2_X1 U393 ( .A1(n638), .A2(n592), .ZN(n427) );
  XNOR2_X1 U394 ( .A(n393), .B(n392), .ZN(n754) );
  XOR2_X1 U395 ( .A(n559), .B(n558), .Z(n598) );
  OR2_X1 U396 ( .A1(n720), .A2(G902), .ZN(n524) );
  XNOR2_X1 U397 ( .A(n720), .B(n719), .ZN(n721) );
  OR2_X1 U398 ( .A1(n750), .A2(n749), .ZN(n393) );
  XNOR2_X1 U399 ( .A(n375), .B(n540), .ZN(n583) );
  NAND2_X1 U400 ( .A1(n389), .A2(n372), .ZN(n357) );
  NAND2_X1 U401 ( .A1(n389), .A2(n372), .ZN(n801) );
  XNOR2_X2 U402 ( .A(n529), .B(n370), .ZN(n432) );
  XNOR2_X2 U403 ( .A(n432), .B(n528), .ZN(n712) );
  XNOR2_X2 U404 ( .A(n435), .B(n516), .ZN(n528) );
  BUF_X1 U405 ( .A(n529), .Z(n358) );
  NOR2_X1 U406 ( .A1(n676), .A2(n675), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n594), .B(n584), .ZN(n360) );
  BUF_X1 U408 ( .A(n594), .Z(n361) );
  XNOR2_X1 U409 ( .A(n594), .B(n584), .ZN(n620) );
  AND2_X1 U410 ( .A1(n658), .A2(n657), .ZN(n699) );
  XNOR2_X2 U411 ( .A(n800), .B(G146), .ZN(n522) );
  XNOR2_X2 U412 ( .A(n464), .B(n535), .ZN(n800) );
  NAND2_X1 U413 ( .A1(n449), .A2(n448), .ZN(n658) );
  NAND2_X1 U414 ( .A1(n462), .A2(n461), .ZN(n457) );
  XOR2_X1 U415 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n545) );
  INV_X1 U416 ( .A(G134), .ZN(n501) );
  XNOR2_X1 U417 ( .A(n680), .B(KEYINPUT45), .ZN(n681) );
  XNOR2_X1 U418 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n621) );
  INV_X1 U419 ( .A(n621), .ZN(n451) );
  INV_X1 U420 ( .A(n448), .ZN(n442) );
  XNOR2_X1 U421 ( .A(G902), .B(KEYINPUT90), .ZN(n409) );
  INV_X1 U422 ( .A(KEYINPUT8), .ZN(n489) );
  INV_X1 U423 ( .A(KEYINPUT113), .ZN(n392) );
  INV_X1 U424 ( .A(KEYINPUT1), .ZN(n411) );
  INV_X1 U425 ( .A(G902), .ZN(n615) );
  XNOR2_X1 U426 ( .A(G119), .B(G116), .ZN(n516) );
  XNOR2_X1 U427 ( .A(n517), .B(KEYINPUT3), .ZN(n435) );
  XNOR2_X1 U428 ( .A(G119), .B(G128), .ZN(n486) );
  NOR2_X1 U429 ( .A1(n660), .A2(n670), .ZN(n423) );
  XNOR2_X1 U430 ( .A(n796), .B(KEYINPUT85), .ZN(n607) );
  XOR2_X1 U431 ( .A(G122), .B(G104), .Z(n552) );
  XNOR2_X1 U432 ( .A(G113), .B(G143), .ZN(n551) );
  XNOR2_X1 U433 ( .A(n546), .B(n429), .ZN(n550) );
  XNOR2_X1 U434 ( .A(KEYINPUT101), .B(KEYINPUT11), .ZN(n544) );
  XNOR2_X1 U435 ( .A(n547), .B(n465), .ZN(n464) );
  XNOR2_X1 U436 ( .A(n499), .B(n501), .ZN(n465) );
  INV_X1 U437 ( .A(G137), .ZN(n499) );
  INV_X1 U438 ( .A(KEYINPUT2), .ZN(n479) );
  XNOR2_X1 U439 ( .A(n566), .B(KEYINPUT4), .ZN(n535) );
  NAND2_X1 U440 ( .A1(n397), .A2(n367), .ZN(n394) );
  INV_X1 U441 ( .A(n681), .ZN(n413) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n507) );
  INV_X1 U443 ( .A(KEYINPUT75), .ZN(n379) );
  INV_X1 U444 ( .A(KEYINPUT76), .ZN(n469) );
  OR2_X2 U445 ( .A1(n620), .A2(n371), .ZN(n448) );
  OR2_X1 U446 ( .A1(n363), .A2(n451), .ZN(n450) );
  XOR2_X1 U447 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n480) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n548) );
  XNOR2_X1 U449 ( .A(KEYINPUT104), .B(KEYINPUT7), .ZN(n562) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n515), .B(KEYINPUT93), .ZN(n749) );
  NOR2_X1 U452 ( .A1(n754), .A2(n753), .ZN(n391) );
  OR2_X1 U453 ( .A1(n588), .A2(n628), .ZN(n406) );
  XNOR2_X1 U454 ( .A(n408), .B(KEYINPUT97), .ZN(n656) );
  XOR2_X1 U455 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n491) );
  XNOR2_X1 U456 ( .A(n730), .B(KEYINPUT59), .ZN(n731) );
  INV_X1 U457 ( .A(KEYINPUT109), .ZN(n436) );
  INV_X1 U458 ( .A(KEYINPUT56), .ZN(n430) );
  AND2_X1 U459 ( .A1(n406), .A2(n629), .ZN(n362) );
  OR2_X1 U460 ( .A1(n619), .A2(n618), .ZN(n363) );
  INV_X1 U461 ( .A(n717), .ZN(n388) );
  XNOR2_X1 U462 ( .A(G143), .B(G128), .ZN(n566) );
  XOR2_X1 U463 ( .A(n726), .B(n725), .Z(n364) );
  AND2_X1 U464 ( .A1(n460), .A2(n659), .ZN(n365) );
  AND2_X1 U465 ( .A1(n587), .A2(n586), .ZN(n366) );
  AND2_X1 U466 ( .A1(n415), .A2(n413), .ZN(n367) );
  AND2_X1 U467 ( .A1(n668), .A2(n667), .ZN(n368) );
  AND2_X1 U468 ( .A1(n471), .A2(G210), .ZN(n369) );
  XOR2_X1 U469 ( .A(KEYINPUT16), .B(G122), .Z(n370) );
  NAND2_X1 U470 ( .A1(n363), .A2(n451), .ZN(n371) );
  BUF_X1 U471 ( .A(n644), .Z(n588) );
  AND2_X1 U472 ( .A1(n388), .A2(n798), .ZN(n372) );
  XNOR2_X1 U473 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n373) );
  XOR2_X1 U474 ( .A(n381), .B(n436), .Z(n374) );
  INV_X1 U475 ( .A(KEYINPUT34), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n409), .B(KEYINPUT15), .ZN(n682) );
  NOR2_X2 U477 ( .A1(n583), .A2(n749), .ZN(n384) );
  OR2_X2 U478 ( .A1(n687), .A2(n376), .ZN(n375) );
  INV_X1 U479 ( .A(n682), .ZN(n376) );
  XNOR2_X1 U480 ( .A(n470), .B(n469), .ZN(n527) );
  NAND2_X1 U481 ( .A1(n656), .A2(n513), .ZN(n470) );
  NOR2_X1 U482 ( .A1(n608), .A2(n366), .ZN(n468) );
  NAND2_X1 U483 ( .A1(n395), .A2(n394), .ZN(n377) );
  BUF_X1 U484 ( .A(n472), .Z(n378) );
  NAND2_X1 U485 ( .A1(n395), .A2(n394), .ZN(n706) );
  AND2_X1 U486 ( .A1(n414), .A2(n359), .ZN(n397) );
  NAND2_X1 U487 ( .A1(n679), .A2(n678), .ZN(n414) );
  NAND2_X1 U488 ( .A1(n404), .A2(n403), .ZN(n381) );
  NAND2_X1 U489 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X2 U490 ( .A1(n443), .A2(n438), .ZN(n383) );
  NAND2_X1 U491 ( .A1(n443), .A2(n438), .ZN(n475) );
  XNOR2_X1 U492 ( .A(n402), .B(n436), .ZN(n635) );
  XNOR2_X2 U493 ( .A(n424), .B(KEYINPUT106), .ZN(n665) );
  XNOR2_X1 U494 ( .A(n647), .B(n646), .ZN(n382) );
  XNOR2_X1 U495 ( .A(n647), .B(n646), .ZN(n748) );
  NOR2_X1 U496 ( .A1(n738), .A2(G902), .ZN(n505) );
  BUF_X1 U497 ( .A(n706), .Z(n426) );
  AND2_X1 U498 ( .A1(n389), .A2(n388), .ZN(n685) );
  NOR2_X2 U499 ( .A1(n597), .A2(n588), .ZN(n796) );
  XNOR2_X2 U500 ( .A(n384), .B(KEYINPUT89), .ZN(n594) );
  NAND2_X1 U501 ( .A1(n405), .A2(KEYINPUT108), .ZN(n403) );
  NAND2_X1 U502 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U503 ( .A1(n665), .A2(n368), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n425), .A2(n385), .ZN(n676) );
  AND2_X1 U505 ( .A1(n638), .A2(n631), .ZN(n474) );
  AND2_X2 U506 ( .A1(n386), .A2(n446), .ZN(n443) );
  NAND2_X1 U507 ( .A1(n445), .A2(n444), .ZN(n386) );
  NAND2_X1 U508 ( .A1(n458), .A2(n457), .ZN(n668) );
  XNOR2_X2 U509 ( .A(n387), .B(n373), .ZN(n793) );
  NAND2_X1 U510 ( .A1(n658), .A2(n654), .ZN(n387) );
  XNOR2_X2 U511 ( .A(n466), .B(n390), .ZN(n389) );
  AND2_X2 U512 ( .A1(n396), .A2(n398), .ZN(n395) );
  NAND2_X1 U513 ( .A1(n400), .A2(n681), .ZN(n396) );
  NAND2_X1 U514 ( .A1(n399), .A2(n681), .ZN(n398) );
  INV_X1 U515 ( .A(n428), .ZN(n399) );
  NAND2_X1 U516 ( .A1(n414), .A2(n415), .ZN(n400) );
  AND2_X2 U517 ( .A1(n401), .A2(n362), .ZN(n404) );
  NAND2_X1 U518 ( .A1(n383), .A2(n407), .ZN(n401) );
  INV_X1 U519 ( .A(n383), .ZN(n405) );
  AND2_X1 U520 ( .A1(n588), .A2(n628), .ZN(n407) );
  NAND2_X1 U521 ( .A1(n410), .A2(n577), .ZN(n408) );
  INV_X1 U522 ( .A(n760), .ZN(n410) );
  XNOR2_X1 U523 ( .A(n577), .B(n411), .ZN(n644) );
  XNOR2_X2 U524 ( .A(n505), .B(n412), .ZN(n577) );
  INV_X1 U525 ( .A(G469), .ZN(n412) );
  NAND2_X1 U526 ( .A1(n664), .A2(n677), .ZN(n415) );
  NOR2_X1 U527 ( .A1(n748), .A2(n420), .ZN(n418) );
  OR2_X1 U528 ( .A1(n658), .A2(n422), .ZN(n419) );
  NAND2_X1 U529 ( .A1(n416), .A2(n421), .ZN(n652) );
  NOR2_X1 U530 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U531 ( .A1(n419), .A2(n649), .ZN(n417) );
  NAND2_X1 U532 ( .A1(n658), .A2(n422), .ZN(n420) );
  NAND2_X1 U533 ( .A1(n382), .A2(KEYINPUT34), .ZN(n421) );
  NAND2_X1 U534 ( .A1(n423), .A2(n665), .ZN(n663) );
  INV_X1 U535 ( .A(n449), .ZN(n445) );
  NAND2_X1 U536 ( .A1(n643), .A2(n642), .ZN(n424) );
  NOR2_X2 U537 ( .A1(n426), .A2(n686), .ZN(n746) );
  AND2_X2 U538 ( .A1(n472), .A2(n471), .ZN(n737) );
  NAND2_X1 U539 ( .A1(n745), .A2(n376), .ZN(n453) );
  NAND2_X1 U540 ( .A1(n653), .A2(n645), .ZN(n647) );
  INV_X1 U541 ( .A(n547), .ZN(n429) );
  XNOR2_X1 U542 ( .A(n431), .B(n430), .ZN(G51) );
  NAND2_X1 U543 ( .A1(n693), .A2(n733), .ZN(n431) );
  NAND2_X1 U544 ( .A1(n378), .A2(n369), .ZN(n691) );
  NAND2_X1 U545 ( .A1(n737), .A2(G472), .ZN(n722) );
  NAND2_X1 U546 ( .A1(n737), .A2(G475), .ZN(n732) );
  XNOR2_X2 U547 ( .A(n434), .B(n433), .ZN(n529) );
  XNOR2_X2 U548 ( .A(G110), .B(G107), .ZN(n433) );
  XNOR2_X2 U549 ( .A(G104), .B(G101), .ZN(n434) );
  AND2_X2 U550 ( .A1(n437), .A2(n450), .ZN(n449) );
  NAND2_X1 U551 ( .A1(n360), .A2(n621), .ZN(n437) );
  NAND2_X1 U552 ( .A1(n442), .A2(n444), .ZN(n441) );
  NAND2_X1 U553 ( .A1(n440), .A2(n476), .ZN(n439) );
  INV_X1 U554 ( .A(n625), .ZN(n440) );
  NAND2_X1 U555 ( .A1(n447), .A2(n449), .ZN(n446) );
  AND2_X2 U556 ( .A1(n448), .A2(n476), .ZN(n447) );
  NAND2_X1 U557 ( .A1(n454), .A2(n452), .ZN(n472) );
  NAND2_X1 U558 ( .A1(n453), .A2(n473), .ZN(n452) );
  NOR2_X2 U559 ( .A1(n377), .A2(n357), .ZN(n745) );
  NAND2_X1 U560 ( .A1(n455), .A2(n376), .ZN(n454) );
  NAND2_X1 U561 ( .A1(n456), .A2(n479), .ZN(n455) );
  NAND2_X1 U562 ( .A1(n477), .A2(n478), .ZN(n456) );
  NAND2_X1 U563 ( .A1(n793), .A2(KEYINPUT99), .ZN(n459) );
  NAND2_X1 U564 ( .A1(n699), .A2(KEYINPUT99), .ZN(n460) );
  NOR2_X1 U565 ( .A1(n699), .A2(KEYINPUT99), .ZN(n461) );
  INV_X1 U566 ( .A(n793), .ZN(n462) );
  XNOR2_X2 U567 ( .A(G125), .B(G146), .ZN(n531) );
  NAND2_X1 U568 ( .A1(n463), .A2(n792), .ZN(n798) );
  XNOR2_X1 U569 ( .A(n543), .B(n542), .ZN(n463) );
  NAND2_X1 U570 ( .A1(n468), .A2(n467), .ZN(n466) );
  XNOR2_X1 U571 ( .A(n582), .B(KEYINPUT46), .ZN(n467) );
  INV_X1 U572 ( .A(n746), .ZN(n471) );
  INV_X1 U573 ( .A(KEYINPUT84), .ZN(n473) );
  NAND2_X1 U574 ( .A1(n475), .A2(n638), .ZN(n640) );
  NAND2_X1 U575 ( .A1(n474), .A2(n383), .ZN(n633) );
  INV_X1 U576 ( .A(n627), .ZN(n476) );
  INV_X1 U577 ( .A(n706), .ZN(n477) );
  NOR2_X1 U578 ( .A1(n602), .A2(n750), .ZN(n543) );
  NAND2_X1 U579 ( .A1(n682), .A2(G234), .ZN(n481) );
  XNOR2_X1 U580 ( .A(n481), .B(n480), .ZN(n495) );
  NAND2_X1 U581 ( .A1(n495), .A2(G221), .ZN(n483) );
  INV_X1 U582 ( .A(KEYINPUT21), .ZN(n482) );
  XNOR2_X1 U583 ( .A(n483), .B(n482), .ZN(n764) );
  INV_X1 U584 ( .A(KEYINPUT96), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n764), .B(n484), .ZN(n622) );
  XNOR2_X1 U586 ( .A(G140), .B(KEYINPUT10), .ZN(n485) );
  XNOR2_X1 U587 ( .A(n531), .B(n485), .ZN(n799) );
  XOR2_X1 U588 ( .A(G110), .B(G137), .Z(n487) );
  XNOR2_X1 U589 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U590 ( .A(n799), .B(n488), .ZN(n494) );
  NAND2_X1 U591 ( .A1(n805), .A2(G234), .ZN(n490) );
  XNOR2_X1 U592 ( .A(n490), .B(n489), .ZN(n565) );
  AND2_X1 U593 ( .A1(n565), .A2(G221), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n494), .B(n493), .ZN(n726) );
  NAND2_X1 U596 ( .A1(n726), .A2(n615), .ZN(n498) );
  NAND2_X1 U597 ( .A1(n495), .A2(G217), .ZN(n496) );
  XNOR2_X1 U598 ( .A(n496), .B(KEYINPUT25), .ZN(n497) );
  XNOR2_X2 U599 ( .A(n498), .B(n497), .ZN(n762) );
  OR2_X1 U600 ( .A1(n622), .A2(n762), .ZN(n760) );
  XNOR2_X2 U601 ( .A(G131), .B(KEYINPUT70), .ZN(n500) );
  NAND2_X1 U602 ( .A1(n805), .A2(G227), .ZN(n502) );
  XNOR2_X1 U603 ( .A(n502), .B(G140), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n358), .B(n503), .ZN(n504) );
  XNOR2_X1 U605 ( .A(n522), .B(n504), .ZN(n738) );
  INV_X1 U606 ( .A(KEYINPUT14), .ZN(n506) );
  XNOR2_X1 U607 ( .A(n507), .B(n506), .ZN(n616) );
  INV_X1 U608 ( .A(G952), .ZN(n692) );
  OR2_X1 U609 ( .A1(n616), .A2(n692), .ZN(n777) );
  NOR2_X1 U610 ( .A1(n777), .A2(G953), .ZN(n619) );
  NAND2_X1 U611 ( .A1(G953), .A2(G902), .ZN(n508) );
  NOR2_X1 U612 ( .A1(n616), .A2(n508), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n509), .B(KEYINPUT111), .ZN(n510) );
  NOR2_X1 U614 ( .A1(G900), .A2(n510), .ZN(n511) );
  NOR2_X1 U615 ( .A1(n619), .A2(n511), .ZN(n512) );
  XNOR2_X1 U616 ( .A(n512), .B(KEYINPUT80), .ZN(n573) );
  INV_X1 U617 ( .A(n573), .ZN(n513) );
  INV_X1 U618 ( .A(G237), .ZN(n514) );
  NAND2_X1 U619 ( .A1(n615), .A2(n514), .ZN(n538) );
  NAND2_X1 U620 ( .A1(n538), .A2(G214), .ZN(n515) );
  XNOR2_X2 U621 ( .A(G113), .B(KEYINPUT72), .ZN(n517) );
  XOR2_X1 U622 ( .A(G101), .B(KEYINPUT5), .Z(n519) );
  NAND2_X1 U623 ( .A1(n548), .A2(G210), .ZN(n518) );
  XNOR2_X1 U624 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U625 ( .A(n528), .B(n520), .ZN(n521) );
  XNOR2_X1 U626 ( .A(n522), .B(n521), .ZN(n720) );
  XNOR2_X1 U627 ( .A(KEYINPUT73), .B(G472), .ZN(n523) );
  XNOR2_X2 U628 ( .A(n524), .B(n523), .ZN(n655) );
  NOR2_X1 U629 ( .A1(n749), .A2(n655), .ZN(n525) );
  XNOR2_X1 U630 ( .A(KEYINPUT30), .B(n525), .ZN(n526) );
  NAND2_X1 U631 ( .A1(n527), .A2(n526), .ZN(n602) );
  XNOR2_X1 U632 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n530) );
  XNOR2_X1 U633 ( .A(n531), .B(n530), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n805), .A2(G224), .ZN(n532) );
  XNOR2_X1 U635 ( .A(n532), .B(KEYINPUT91), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n534), .B(n533), .ZN(n536) );
  XNOR2_X1 U637 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U638 ( .A(n712), .B(n537), .ZN(n687) );
  NAND2_X1 U639 ( .A1(n538), .A2(G210), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n539), .B(KEYINPUT92), .ZN(n540) );
  BUF_X1 U641 ( .A(n583), .Z(n541) );
  XOR2_X1 U642 ( .A(KEYINPUT38), .B(n541), .Z(n750) );
  INV_X1 U643 ( .A(KEYINPUT39), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U645 ( .A1(G214), .A2(n548), .ZN(n549) );
  XNOR2_X1 U646 ( .A(n550), .B(n549), .ZN(n555) );
  XNOR2_X1 U647 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U648 ( .A(n799), .B(n553), .ZN(n554) );
  XNOR2_X1 U649 ( .A(n555), .B(n554), .ZN(n730) );
  NOR2_X1 U650 ( .A1(n730), .A2(G902), .ZN(n559) );
  XOR2_X1 U651 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n557) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(G475), .ZN(n556) );
  XNOR2_X1 U653 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U654 ( .A(G122), .B(G107), .Z(n561) );
  XNOR2_X1 U655 ( .A(G116), .B(G134), .ZN(n560) );
  XNOR2_X1 U656 ( .A(n561), .B(n560), .ZN(n564) );
  XNOR2_X1 U657 ( .A(n562), .B(KEYINPUT9), .ZN(n563) );
  XNOR2_X1 U658 ( .A(n564), .B(n563), .ZN(n570) );
  NAND2_X1 U659 ( .A1(n565), .A2(G217), .ZN(n568) );
  INV_X1 U660 ( .A(n566), .ZN(n567) );
  XNOR2_X1 U661 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U662 ( .A(n570), .B(n569), .ZN(n727) );
  NOR2_X1 U663 ( .A1(G902), .A2(n727), .ZN(n571) );
  XOR2_X1 U664 ( .A(G478), .B(n571), .Z(n599) );
  NOR2_X1 U665 ( .A1(n598), .A2(n599), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n572), .B(KEYINPUT40), .ZN(n812) );
  NAND2_X1 U667 ( .A1(n762), .A2(n764), .ZN(n574) );
  NOR2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n575), .B(KEYINPUT71), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n655), .A2(n592), .ZN(n576) );
  XNOR2_X1 U671 ( .A(KEYINPUT28), .B(n576), .ZN(n578) );
  NAND2_X1 U672 ( .A1(n578), .A2(n577), .ZN(n585) );
  INV_X1 U673 ( .A(n599), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n598), .A2(n579), .ZN(n580) );
  XNOR2_X1 U675 ( .A(n580), .B(KEYINPUT105), .ZN(n624) );
  INV_X1 U676 ( .A(n624), .ZN(n753) );
  NOR2_X1 U677 ( .A1(n585), .A2(n779), .ZN(n581) );
  XNOR2_X1 U678 ( .A(n581), .B(KEYINPUT42), .ZN(n811) );
  NOR2_X1 U679 ( .A1(n812), .A2(n811), .ZN(n582) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n584) );
  NOR2_X1 U681 ( .A1(n585), .A2(n360), .ZN(n790) );
  XOR2_X1 U682 ( .A(KEYINPUT47), .B(n790), .Z(n587) );
  AND2_X1 U683 ( .A1(n598), .A2(n599), .ZN(n792) );
  NOR2_X1 U684 ( .A1(n590), .A2(n792), .ZN(n755) );
  NAND2_X1 U685 ( .A1(n790), .A2(n755), .ZN(n586) );
  INV_X1 U686 ( .A(KEYINPUT110), .ZN(n589) );
  XNOR2_X1 U687 ( .A(n590), .B(n589), .ZN(n694) );
  INV_X1 U688 ( .A(KEYINPUT6), .ZN(n591) );
  XNOR2_X1 U689 ( .A(n655), .B(n591), .ZN(n638) );
  NOR2_X2 U690 ( .A1(n694), .A2(n593), .ZN(n609) );
  INV_X1 U691 ( .A(n361), .ZN(n595) );
  NAND2_X1 U692 ( .A1(n609), .A2(n595), .ZN(n596) );
  XNOR2_X1 U693 ( .A(n596), .B(KEYINPUT36), .ZN(n597) );
  INV_X1 U694 ( .A(n598), .ZN(n600) );
  NAND2_X1 U695 ( .A1(n600), .A2(n599), .ZN(n648) );
  OR2_X1 U696 ( .A1(n648), .A2(n541), .ZN(n601) );
  NOR2_X1 U697 ( .A1(n602), .A2(n601), .ZN(n696) );
  XNOR2_X1 U698 ( .A(n696), .B(KEYINPUT83), .ZN(n604) );
  NAND2_X1 U699 ( .A1(KEYINPUT47), .A2(n755), .ZN(n603) );
  NAND2_X1 U700 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U701 ( .A(KEYINPUT82), .B(n605), .Z(n606) );
  NAND2_X1 U702 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U703 ( .A1(n588), .A2(n609), .ZN(n610) );
  NOR2_X1 U704 ( .A1(n749), .A2(n610), .ZN(n611) );
  XNOR2_X1 U705 ( .A(n611), .B(KEYINPUT43), .ZN(n613) );
  INV_X1 U706 ( .A(n541), .ZN(n612) );
  NOR2_X1 U707 ( .A1(n613), .A2(n612), .ZN(n717) );
  INV_X1 U708 ( .A(G898), .ZN(n708) );
  NAND2_X1 U709 ( .A1(n708), .A2(G953), .ZN(n614) );
  XNOR2_X1 U710 ( .A(n614), .B(KEYINPUT94), .ZN(n713) );
  OR2_X1 U711 ( .A1(n713), .A2(n615), .ZN(n617) );
  NOR2_X1 U712 ( .A1(n617), .A2(n616), .ZN(n618) );
  INV_X1 U713 ( .A(n622), .ZN(n623) );
  AND2_X1 U714 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U715 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n626) );
  XNOR2_X1 U716 ( .A(n626), .B(KEYINPUT66), .ZN(n627) );
  INV_X1 U717 ( .A(n588), .ZN(n641) );
  INV_X1 U718 ( .A(KEYINPUT108), .ZN(n628) );
  AND2_X1 U719 ( .A1(n655), .A2(n762), .ZN(n629) );
  NAND2_X1 U720 ( .A1(n762), .A2(n641), .ZN(n630) );
  XNOR2_X1 U721 ( .A(n630), .B(KEYINPUT107), .ZN(n631) );
  XNOR2_X1 U722 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n632) );
  INV_X1 U723 ( .A(n705), .ZN(n634) );
  INV_X1 U724 ( .A(KEYINPUT88), .ZN(n636) );
  XNOR2_X2 U725 ( .A(n637), .B(n636), .ZN(n677) );
  INV_X1 U726 ( .A(n638), .ZN(n645) );
  INV_X1 U727 ( .A(KEYINPUT86), .ZN(n639) );
  XNOR2_X1 U728 ( .A(n640), .B(n639), .ZN(n643) );
  NOR2_X1 U729 ( .A1(n762), .A2(n641), .ZN(n642) );
  INV_X1 U730 ( .A(KEYINPUT33), .ZN(n646) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT79), .ZN(n649) );
  INV_X1 U732 ( .A(KEYINPUT78), .ZN(n650) );
  XNOR2_X1 U733 ( .A(n650), .B(KEYINPUT35), .ZN(n651) );
  XNOR2_X2 U734 ( .A(n652), .B(n651), .ZN(n718) );
  NAND2_X1 U735 ( .A1(n718), .A2(KEYINPUT87), .ZN(n660) );
  INV_X1 U736 ( .A(n655), .ZN(n767) );
  NAND2_X1 U737 ( .A1(n767), .A2(n653), .ZN(n770) );
  INV_X1 U738 ( .A(n770), .ZN(n654) );
  AND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n657) );
  INV_X1 U740 ( .A(n755), .ZN(n659) );
  INV_X1 U741 ( .A(n668), .ZN(n670) );
  INV_X1 U742 ( .A(KEYINPUT44), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n718), .A2(n666), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(KEYINPUT68), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n664) );
  INV_X1 U746 ( .A(n665), .ZN(n674) );
  AND2_X1 U747 ( .A1(n666), .A2(KEYINPUT87), .ZN(n667) );
  INV_X1 U748 ( .A(n718), .ZN(n669) );
  INV_X1 U749 ( .A(KEYINPUT87), .ZN(n673) );
  AND2_X1 U750 ( .A1(n673), .A2(KEYINPUT44), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n669), .A2(n678), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n670), .A2(n673), .ZN(n671) );
  INV_X1 U753 ( .A(n677), .ZN(n679) );
  INV_X1 U754 ( .A(KEYINPUT64), .ZN(n680) );
  NAND2_X1 U755 ( .A1(n798), .A2(KEYINPUT2), .ZN(n683) );
  XNOR2_X1 U756 ( .A(n683), .B(KEYINPUT81), .ZN(n684) );
  NAND2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n686) );
  BUF_X1 U758 ( .A(n687), .Z(n689) );
  XNOR2_X1 U759 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n688) );
  XNOR2_X1 U760 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n692), .A2(G953), .ZN(n733) );
  INV_X1 U763 ( .A(n694), .ZN(n789) );
  NAND2_X1 U764 ( .A1(n699), .A2(n789), .ZN(n695) );
  XNOR2_X1 U765 ( .A(n695), .B(G104), .ZN(G6) );
  XOR2_X1 U766 ( .A(G143), .B(n696), .Z(G45) );
  XOR2_X1 U767 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n698) );
  XNOR2_X1 U768 ( .A(G107), .B(KEYINPUT27), .ZN(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n701) );
  NAND2_X1 U770 ( .A1(n699), .A2(n792), .ZN(n700) );
  XOR2_X1 U771 ( .A(n701), .B(n700), .Z(G9) );
  XNOR2_X1 U772 ( .A(G113), .B(KEYINPUT117), .ZN(n703) );
  NAND2_X1 U773 ( .A1(n793), .A2(n789), .ZN(n702) );
  XOR2_X1 U774 ( .A(n703), .B(n702), .Z(G15) );
  XNOR2_X1 U775 ( .A(G119), .B(KEYINPUT125), .ZN(n704) );
  XNOR2_X1 U776 ( .A(n705), .B(n704), .ZN(G21) );
  NOR2_X1 U777 ( .A1(n426), .A2(G953), .ZN(n711) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n707) );
  XOR2_X1 U779 ( .A(n707), .B(KEYINPUT61), .Z(n709) );
  NOR2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n716) );
  XOR2_X1 U782 ( .A(KEYINPUT123), .B(n712), .Z(n714) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U784 ( .A(n716), .B(n715), .ZN(G69) );
  XNOR2_X1 U785 ( .A(n665), .B(G101), .ZN(G3) );
  XOR2_X1 U786 ( .A(G140), .B(n717), .Z(G42) );
  XOR2_X1 U787 ( .A(n374), .B(G110), .Z(G12) );
  XNOR2_X1 U788 ( .A(n718), .B(G122), .ZN(G24) );
  XOR2_X1 U789 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n719) );
  XNOR2_X1 U790 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U791 ( .A1(n723), .A2(n733), .ZN(n724) );
  XNOR2_X1 U792 ( .A(n724), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U793 ( .A1(n737), .A2(G217), .ZN(n725) );
  INV_X1 U794 ( .A(n733), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n364), .A2(n743), .ZN(G66) );
  NAND2_X1 U796 ( .A1(n356), .A2(G478), .ZN(n728) );
  XNOR2_X1 U797 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U798 ( .A1(n729), .A2(n743), .ZN(G63) );
  XNOR2_X1 U799 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U800 ( .A1(n734), .A2(n733), .ZN(n736) );
  XOR2_X1 U801 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n735) );
  XNOR2_X1 U802 ( .A(n736), .B(n735), .ZN(G60) );
  NAND2_X1 U803 ( .A1(n356), .A2(G469), .ZN(n742) );
  XNOR2_X1 U804 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n739) );
  XNOR2_X1 U805 ( .A(n739), .B(KEYINPUT58), .ZN(n740) );
  XNOR2_X1 U806 ( .A(n738), .B(n740), .ZN(n741) );
  XNOR2_X1 U807 ( .A(n742), .B(n741), .ZN(n744) );
  NOR2_X1 U808 ( .A1(n744), .A2(n743), .ZN(G54) );
  NOR2_X1 U809 ( .A1(n745), .A2(KEYINPUT2), .ZN(n747) );
  NOR2_X1 U810 ( .A1(n747), .A2(n746), .ZN(n784) );
  NAND2_X1 U811 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U812 ( .A(KEYINPUT119), .B(n751), .ZN(n752) );
  NOR2_X1 U813 ( .A1(n753), .A2(n752), .ZN(n757) );
  NOR2_X1 U814 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U815 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U816 ( .A(n758), .B(KEYINPUT120), .ZN(n759) );
  NOR2_X1 U817 ( .A1(n382), .A2(n759), .ZN(n775) );
  NAND2_X1 U818 ( .A1(n588), .A2(n760), .ZN(n761) );
  XNOR2_X1 U819 ( .A(n761), .B(KEYINPUT50), .ZN(n769) );
  INV_X1 U820 ( .A(n762), .ZN(n763) );
  NOR2_X1 U821 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U822 ( .A(KEYINPUT49), .B(n765), .Z(n766) );
  NOR2_X1 U823 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U824 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U825 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U826 ( .A(KEYINPUT51), .B(n772), .ZN(n773) );
  NOR2_X1 U827 ( .A1(n779), .A2(n773), .ZN(n774) );
  NOR2_X1 U828 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U829 ( .A(n776), .B(KEYINPUT52), .ZN(n778) );
  OR2_X1 U830 ( .A1(n778), .A2(n777), .ZN(n782) );
  NOR2_X1 U831 ( .A1(n779), .A2(n382), .ZN(n780) );
  NOR2_X1 U832 ( .A1(n780), .A2(G953), .ZN(n781) );
  NAND2_X1 U833 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U834 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U835 ( .A(n785), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U836 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n787) );
  NAND2_X1 U837 ( .A1(n790), .A2(n792), .ZN(n786) );
  XNOR2_X1 U838 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U839 ( .A(G128), .B(n788), .ZN(G30) );
  NAND2_X1 U840 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U841 ( .A(n791), .B(G146), .ZN(G48) );
  NAND2_X1 U842 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U843 ( .A(n794), .B(KEYINPUT118), .ZN(n795) );
  XNOR2_X1 U844 ( .A(G116), .B(n795), .ZN(G18) );
  XNOR2_X1 U845 ( .A(G125), .B(n796), .ZN(n797) );
  XNOR2_X1 U846 ( .A(n797), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U847 ( .A(G134), .B(n798), .ZN(G36) );
  XNOR2_X1 U848 ( .A(n800), .B(n799), .ZN(n803) );
  XNOR2_X1 U849 ( .A(n803), .B(n357), .ZN(n802) );
  NOR2_X1 U850 ( .A1(G953), .A2(n802), .ZN(n808) );
  XNOR2_X1 U851 ( .A(G227), .B(n803), .ZN(n804) );
  NAND2_X1 U852 ( .A1(n804), .A2(G900), .ZN(n806) );
  NOR2_X1 U853 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U854 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U855 ( .A(KEYINPUT124), .B(n809), .ZN(G72) );
  XOR2_X1 U856 ( .A(G137), .B(KEYINPUT126), .Z(n810) );
  XNOR2_X1 U857 ( .A(n811), .B(n810), .ZN(G39) );
  XNOR2_X1 U858 ( .A(G131), .B(KEYINPUT127), .ZN(n813) );
  XNOR2_X1 U859 ( .A(n813), .B(n812), .ZN(G33) );
endmodule

