//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT64), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n461), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n464), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n461), .A2(new_n465), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(G136), .B2(new_n469), .ZN(G162));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n459), .A2(new_n460), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n465), .ZN(new_n481));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(G102), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT4), .A2(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n461), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n461), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n483), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  XNOR2_X1  g068(.A(KEYINPUT6), .B(G651), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G50), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G651), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n498), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n495), .A2(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(KEYINPUT65), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(KEYINPUT66), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n519), .B1(new_n501), .B2(new_n502), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G63), .ZN(new_n523));
  NAND3_X1  g098(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n497), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n503), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  AND3_X1   g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT67), .B(G51), .Z(new_n529));
  OAI221_X1 g104(.A(new_n527), .B1(KEYINPUT7), .B2(new_n528), .C1(new_n495), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n498), .A2(new_n500), .A3(G52), .A4(G543), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n533), .B(new_n534), .C1(new_n503), .C2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n506), .A2(new_n494), .A3(G90), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n533), .B1(new_n538), .B2(new_n534), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n518), .A2(new_n520), .A3(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n497), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n532), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n534), .B1(new_n503), .B2(new_n535), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT68), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n536), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n541), .A2(new_n542), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(KEYINPUT69), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n544), .A2(new_n550), .ZN(G171));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT70), .B(G81), .Z(new_n553));
  OAI22_X1  g128(.A1(new_n495), .A2(new_n552), .B1(new_n503), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT71), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n556));
  OAI221_X1 g131(.A(new_n556), .B1(new_n503), .B2(new_n553), .C1(new_n552), .C2(new_n495), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n521), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  XNOR2_X1  g145(.A(new_n503), .B(KEYINPUT73), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n494), .A2(G53), .A3(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n506), .A2(G65), .ZN(new_n575));
  AND2_X1   g150(.A1(G78), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(G299));
  AND3_X1   g153(.A1(new_n547), .A2(KEYINPUT69), .A3(new_n549), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT69), .B1(new_n547), .B2(new_n549), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT74), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n544), .B2(new_n550), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n571), .A2(G87), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n522), .A2(G74), .ZN(new_n589));
  INV_X1    g164(.A(new_n495), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n589), .A2(G651), .B1(G49), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n506), .A2(G61), .ZN(new_n593));
  INV_X1    g168(.A(G73), .ZN(new_n594));
  INV_X1    g169(.A(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n590), .B2(G48), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n503), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(G305));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n495), .A2(new_n602), .B1(new_n503), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n518), .A2(new_n520), .A3(G60), .ZN(new_n606));
  INV_X1    g181(.A(G72), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n595), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n497), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n606), .B(KEYINPUT76), .C1(new_n607), .C2(new_n595), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(KEYINPUT77), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT77), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n613), .B2(new_n614), .ZN(G290));
  INV_X1    g190(.A(G301), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n616), .A2(KEYINPUT78), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT78), .B1(new_n616), .B2(new_n617), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G54), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n620), .A2(new_n497), .B1(new_n621), .B2(new_n495), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n600), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n571), .A2(KEYINPUT10), .A3(G92), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n618), .B(new_n619), .C1(G868), .C2(new_n630), .ZN(G284));
  OAI211_X1 g206(.A(new_n618), .B(new_n619), .C1(G868), .C2(new_n630), .ZN(G321));
  NAND2_X1  g207(.A1(G299), .A2(new_n617), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G168), .B2(new_n617), .ZN(G280));
  XNOR2_X1  g209(.A(G280), .B(KEYINPUT80), .ZN(G297));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n630), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n467), .A2(new_n480), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT81), .ZN(new_n646));
  AOI22_X1  g221(.A1(G123), .A2(new_n473), .B1(new_n469), .B2(G135), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n648), .A2(new_n465), .A3(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n465), .B2(G111), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n646), .B(new_n654), .C1(G2100), .C2(new_n644), .ZN(G156));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(G14), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT17), .Z(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(new_n673), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n678), .C1(new_n676), .C2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n673), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT18), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n653), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n685), .A2(G2100), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(G2100), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n693), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  AOI211_X1 g272(.A(new_n695), .B(new_n697), .C1(new_n690), .C2(new_n694), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT83), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n588), .A2(new_n591), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT33), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(new_n708), .C1(new_n709), .C2(new_n707), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G1976), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n711), .A2(G1976), .A3(new_n713), .ZN(new_n717));
  MUX2_X1   g292(.A(G6), .B(G305), .S(G16), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT32), .B(G1981), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n707), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n707), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G1971), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(G1971), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n716), .A2(new_n717), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n716), .A2(new_n728), .A3(new_n717), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n608), .A2(new_n609), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n730), .A2(G651), .A3(new_n611), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT77), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n604), .B1(new_n733), .B2(new_n612), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G16), .B2(G24), .ZN(new_n736));
  INV_X1    g311(.A(G1986), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT84), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT84), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n469), .A2(G131), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n473), .A2(G119), .ZN(new_n747));
  OR2_X1    g322(.A1(G95), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n744), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n738), .A2(new_n739), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n727), .A2(new_n729), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT36), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n727), .A2(new_n759), .A3(new_n729), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n743), .A2(G26), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT87), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n469), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n473), .A2(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT86), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n740), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n467), .A2(G105), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT90), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n469), .A2(G141), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n473), .A2(G129), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n707), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT97), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT23), .ZN(new_n791));
  INV_X1    g366(.A(G299), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n707), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1956), .Z(new_n794));
  NAND3_X1  g369(.A1(new_n773), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n564), .A2(new_n707), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n707), .B2(G19), .ZN(new_n797));
  INV_X1    g372(.A(G1341), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n707), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n707), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(G1966), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n797), .B2(new_n798), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n744), .A2(G35), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n744), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n743), .A2(G27), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT95), .Z(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n492), .B2(new_n744), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT96), .B(G2078), .Z(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(G28), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT30), .ZN(new_n816));
  AOI21_X1  g391(.A(G29), .B1(new_n815), .B2(KEYINPUT30), .ZN(new_n817));
  OR2_X1    g392(.A1(KEYINPUT31), .A2(G11), .ZN(new_n818));
  NAND2_X1  g393(.A1(KEYINPUT31), .A2(G11), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n816), .A2(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n652), .B2(new_n743), .ZN(new_n821));
  INV_X1    g396(.A(G2084), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT24), .B(G34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n743), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT88), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n471), .B2(new_n740), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n821), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n813), .A2(new_n814), .A3(new_n827), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n795), .A2(new_n804), .A3(new_n808), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(G115), .A2(G2104), .ZN(new_n830));
  INV_X1    g405(.A(G127), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n461), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G2105), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT25), .Z(new_n835));
  INV_X1    g410(.A(G139), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n835), .C1(new_n836), .C2(new_n481), .ZN(new_n837));
  MUX2_X1   g412(.A(G33), .B(new_n837), .S(G29), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G2072), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT89), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n838), .A2(G2072), .B1(new_n826), .B2(new_n822), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n785), .B2(new_n787), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(KEYINPUT93), .C1(new_n785), .C2(new_n787), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n707), .A2(G5), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G171), .B2(new_n707), .ZN(new_n849));
  INV_X1    g424(.A(G1961), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n801), .A2(G1966), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT94), .Z(new_n853));
  NOR2_X1   g428(.A1(G4), .A2(G16), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT85), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n624), .A2(new_n629), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n707), .ZN(new_n857));
  INV_X1    g432(.A(G1348), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n829), .A2(new_n847), .A3(new_n851), .A4(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT98), .B1(new_n761), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n864));
  AOI211_X1 g439(.A(new_n864), .B(new_n861), .C1(new_n758), .C2(new_n760), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(G311));
  NAND2_X1  g441(.A1(new_n761), .A2(new_n862), .ZN(G150));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n495), .A2(new_n868), .B1(new_n503), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  INV_X1    g446(.A(G67), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n521), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n873), .B2(G651), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n874), .A2(KEYINPUT99), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(KEYINPUT99), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n563), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n564), .A2(new_n874), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n630), .A2(G559), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n883), .A2(new_n884), .A3(G860), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n875), .A2(new_n876), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G860), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT37), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n885), .A2(new_n888), .ZN(G145));
  XNOR2_X1  g464(.A(new_n492), .B(new_n769), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n783), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n837), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n469), .A2(G142), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n473), .A2(G130), .ZN(new_n894));
  NOR2_X1   g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n643), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n751), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT100), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n892), .A2(new_n899), .ZN(new_n903));
  XNOR2_X1  g478(.A(G160), .B(new_n652), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G162), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n903), .B(KEYINPUT101), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n908), .B2(new_n901), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT40), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(G395));
  XNOR2_X1  g487(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n638), .B(KEYINPUT102), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n879), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n856), .A2(new_n792), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n624), .A2(new_n629), .A3(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n624), .A2(new_n629), .A3(G299), .ZN(new_n921));
  AOI21_X1  g496(.A(G299), .B1(new_n624), .B2(new_n629), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n917), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n915), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n913), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n733), .A2(new_n612), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT104), .B1(new_n931), .B2(new_n605), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n933), .B(new_n604), .C1(new_n733), .C2(new_n612), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n709), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G290), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(G288), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(G303), .A2(G305), .ZN(new_n939));
  NAND2_X1  g514(.A1(G303), .A2(G305), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n935), .A2(new_n938), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(KEYINPUT105), .A3(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n935), .B2(new_n938), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n915), .A2(new_n918), .ZN(new_n950));
  INV_X1    g525(.A(new_n913), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n951), .C1(new_n915), .C2(new_n928), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n930), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n930), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n886), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(G868), .B2(new_n956), .ZN(G295));
  OAI21_X1  g532(.A(new_n955), .B1(G868), .B2(new_n956), .ZN(G331));
  XNOR2_X1  g533(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT74), .B1(new_n579), .B2(new_n580), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n544), .A2(new_n582), .A3(new_n550), .ZN(new_n963));
  AOI21_X1  g538(.A(G286), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(G171), .A2(G168), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n879), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(G168), .B1(new_n581), .B2(new_n583), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n877), .A2(new_n878), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n970), .A3(new_n927), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n966), .A2(new_n970), .A3(new_n927), .A4(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n966), .A2(new_n970), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n918), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n948), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n935), .A2(new_n938), .A3(new_n944), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n961), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n971), .A2(new_n972), .B1(new_n975), .B2(new_n918), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n949), .B1(new_n974), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n960), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(KEYINPUT110), .B(new_n960), .C1(new_n981), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n918), .A2(new_n925), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n916), .A2(new_n920), .A3(new_n917), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n966), .A2(new_n970), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n976), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n980), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n982), .A2(new_n949), .A3(new_n974), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n996), .A3(new_n961), .A4(new_n959), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n986), .A2(new_n987), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n981), .A2(new_n983), .A3(new_n960), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n981), .B1(new_n980), .B2(new_n994), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1001), .B(KEYINPUT44), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(G397));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n492), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n464), .A2(new_n468), .A3(G40), .A4(new_n470), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n751), .A2(new_n753), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n750), .A2(new_n754), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n769), .B(G2067), .Z(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1996), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n783), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n776), .A2(G1996), .A3(new_n782), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1015), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n734), .A2(new_n737), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n734), .A2(new_n737), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1012), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT125), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n492), .A2(new_n1028), .A3(new_n1006), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1011), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT117), .B(G1981), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G305), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT118), .B(G86), .Z(new_n1039));
  NAND2_X1  g614(.A1(new_n526), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n700), .B1(new_n597), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT119), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT119), .B(KEYINPUT49), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1036), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n709), .A2(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n715), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1035), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT116), .B1(new_n1031), .B2(G8), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1048), .B(new_n1049), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1036), .B2(new_n1048), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1064), .A2(new_n1030), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1007), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1971), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1029), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1028), .B1(new_n492), .B2(new_n1006), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT50), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G2090), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1030), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1063), .B1(new_n1078), .B2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1027), .A2(new_n1080), .A3(new_n1029), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1011), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1083), .A2(new_n1074), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1062), .ZN(new_n1085));
  OAI21_X1  g660(.A(G8), .B1(new_n1085), .B2(new_n1060), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT115), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1070), .B1(G2090), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1079), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  INV_X1    g671(.A(G2078), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1067), .A2(new_n1097), .A3(new_n1030), .A4(new_n1064), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1090), .A2(new_n850), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1096), .A2(G2078), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1010), .A2(new_n1065), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(G301), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1065), .B(new_n1100), .C1(new_n1104), .C2(KEYINPUT45), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1095), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G171), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1099), .A2(G301), .A3(new_n1105), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(KEYINPUT54), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1056), .A2(new_n1094), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1065), .B1(new_n1104), .B2(KEYINPUT45), .ZN(new_n1113));
  INV_X1    g688(.A(G1966), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1081), .A2(new_n822), .A3(new_n1082), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1113), .A2(new_n1114), .B1(new_n1115), .B2(KEYINPUT120), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1081), .A2(new_n1117), .A3(new_n822), .A4(new_n1082), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(G286), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(KEYINPUT120), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT45), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1064), .A2(new_n1030), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1114), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G168), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(new_n1088), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(new_n1124), .B2(G286), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1026), .B1(new_n1112), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1056), .A2(new_n1094), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1126), .A2(new_n1128), .B1(new_n1130), .B2(new_n1127), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1099), .A2(new_n1105), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1102), .B1(new_n1136), .B2(G301), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1095), .B1(new_n1108), .B2(G171), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1137), .A2(new_n1095), .B1(new_n1138), .B2(new_n1110), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1134), .A2(new_n1135), .A3(KEYINPUT125), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(G1956), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT56), .B(G2072), .Z(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1065), .A2(new_n1067), .A3(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(G299), .B(KEYINPUT57), .Z(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1148), .A2(KEYINPUT61), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1142), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1146), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1153), .A2(new_n1154), .A3(KEYINPUT123), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1149), .B1(new_n1156), .B2(new_n1147), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  AOI21_X1  g733(.A(G1348), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1031), .A2(G2067), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1159), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1159), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1160), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n1166), .A3(KEYINPUT122), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1161), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1164), .A2(new_n1169), .A3(new_n630), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1147), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1148), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT58), .B(G1341), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1031), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(G1996), .B2(new_n1068), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n564), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT59), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1179), .A2(KEYINPUT124), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1177), .B(new_n564), .C1(KEYINPUT124), .C2(new_n1179), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1173), .A2(new_n1174), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(KEYINPUT60), .B(new_n856), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1157), .A2(new_n1170), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1156), .A2(new_n1147), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1162), .A2(new_n1163), .A3(new_n856), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1148), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1133), .A2(new_n1140), .A3(new_n1189), .ZN(new_n1190));
  AOI211_X1 g765(.A(G1976), .B(G288), .C1(new_n1036), .C2(new_n1046), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1191), .A2(new_n1038), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1084), .A2(KEYINPUT115), .A3(new_n1086), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1092), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1195), .B(G8), .C1(new_n1078), .C2(new_n1063), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1193), .A2(new_n1194), .B1(new_n1196), .B2(new_n1125), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1192), .A2(new_n1036), .B1(new_n1197), .B2(new_n1056), .ZN(new_n1198));
  OAI21_X1  g773(.A(G8), .B1(new_n1091), .B2(new_n1063), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1125), .A2(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1036), .A2(new_n1048), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1052), .B(new_n1047), .C1(new_n1201), .C2(new_n1054), .ZN(new_n1202));
  OAI21_X1  g777(.A(KEYINPUT63), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1129), .A2(KEYINPUT62), .A3(new_n1131), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1204), .A2(new_n1134), .A3(new_n1106), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1135), .A2(KEYINPUT62), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1198), .B(new_n1203), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1025), .B1(new_n1190), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT46), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1012), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1209), .B1(new_n1210), .B2(G1996), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1012), .A2(KEYINPUT46), .A3(new_n1018), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1012), .B1(new_n783), .B2(new_n1017), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1214), .B(KEYINPUT47), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1021), .A2(new_n1210), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1210), .A2(new_n1022), .ZN(new_n1217));
  XOR2_X1   g792(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1218));
  AOI21_X1  g793(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1220));
  AOI211_X1 g795(.A(new_n1013), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n769), .A2(G2067), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1012), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1215), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1208), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g800(.A1(new_n907), .A2(new_n909), .ZN(new_n1227));
  NAND4_X1  g801(.A1(new_n686), .A2(new_n671), .A3(G319), .A4(new_n687), .ZN(new_n1228));
  NOR2_X1   g802(.A1(G229), .A2(new_n1228), .ZN(new_n1229));
  AND3_X1   g803(.A1(new_n998), .A2(new_n1227), .A3(new_n1229), .ZN(G308));
  NAND3_X1  g804(.A1(new_n998), .A2(new_n1229), .A3(new_n1227), .ZN(G225));
endmodule


