//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  AOI21_X1  g003(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT18), .A2(G131), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G125), .B(G140), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n201), .B(KEYINPUT76), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n196), .B1(new_n202), .B2(new_n195), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n193), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G113), .B(G122), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n205), .B(G104), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT19), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n194), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n202), .B2(new_n209), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n195), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT74), .B1(new_n201), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT75), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n216), .A2(new_n213), .A3(new_n197), .A4(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n194), .A2(new_n219), .A3(KEYINPUT16), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n218), .A3(G146), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n189), .B2(new_n190), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT86), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G237), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G214), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n188), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT86), .A3(G131), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n191), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n212), .A2(new_n221), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n208), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(G475), .A2(G902), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n238));
  AND4_X1   g052(.A1(new_n238), .A2(new_n224), .A3(new_n231), .A4(new_n233), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT86), .B1(new_n230), .B2(G131), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n223), .B(new_n232), .C1(new_n229), .C2(new_n188), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT17), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n214), .A2(new_n218), .A3(new_n220), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n195), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(new_n221), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n239), .B1(new_n245), .B2(KEYINPUT87), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n242), .A2(new_n247), .A3(new_n244), .A4(new_n221), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n204), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n236), .B(new_n237), .C1(new_n249), .C2(new_n206), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT88), .B1(new_n250), .B2(KEYINPUT20), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n221), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n238), .B1(new_n224), .B2(new_n231), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT87), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n239), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n248), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n204), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n258), .A2(new_n207), .B1(new_n235), .B2(new_n208), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .A4(new_n237), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n250), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n251), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n207), .A2(KEYINPUT89), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n258), .B2(new_n267), .ZN(new_n270));
  OAI21_X1  g084(.A(G475), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT90), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT90), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  XOR2_X1   g089(.A(G128), .B(G143), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT92), .ZN(new_n277));
  XNOR2_X1  g091(.A(G128), .B(G143), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n280), .A3(G134), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n286));
  INV_X1    g100(.A(G122), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(G116), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT91), .A3(G122), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n289), .A2(G122), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT78), .A2(G107), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT78), .A2(G107), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n292), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n299));
  OAI21_X1  g113(.A(G107), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n285), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT13), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n228), .A3(G128), .ZN(new_n303));
  OAI211_X1 g117(.A(G134), .B(new_n303), .C1(new_n276), .C2(new_n302), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n295), .B1(new_n291), .B2(new_n292), .ZN(new_n305));
  INV_X1    g119(.A(new_n296), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n283), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  INV_X1    g122(.A(G217), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n308), .A2(new_n309), .A3(G953), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n301), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n301), .B2(new_n307), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n269), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G478), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT15), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n313), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(G234), .A2(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(G952), .A3(new_n226), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT21), .B(G898), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(G902), .A3(G953), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT93), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n273), .A2(new_n275), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G140), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n226), .A2(G227), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT11), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n282), .B2(G137), .ZN(new_n336));
  INV_X1    g150(.A(G137), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT11), .A3(G134), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n282), .A2(G137), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G131), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n336), .A2(new_n338), .A3(new_n232), .A4(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G101), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n345), .A2(G104), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(new_n295), .B2(G104), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n344), .B(new_n347), .C1(new_n349), .C2(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n195), .A2(G143), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n228), .A2(G146), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT1), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(G128), .ZN(new_n355));
  INV_X1    g169(.A(G128), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n351), .B2(KEYINPUT1), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  INV_X1    g172(.A(G104), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n293), .B2(new_n294), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n344), .B1(new_n360), .B2(new_n346), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n350), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n352), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n228), .C2(G146), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G128), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT64), .B1(new_n351), .B2(KEYINPUT1), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n355), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n350), .B2(new_n362), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n343), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT12), .B1(new_n343), .B2(KEYINPUT81), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n350), .A2(new_n358), .A3(new_n362), .ZN(new_n374));
  OR2_X1    g188(.A1(KEYINPUT78), .A2(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT78), .A2(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(G104), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n348), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT3), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n347), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n361), .B1(new_n381), .B2(new_n344), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n374), .B1(new_n382), .B2(new_n369), .ZN(new_n383));
  INV_X1    g197(.A(new_n372), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n343), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n368), .B2(new_n355), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n374), .A2(new_n387), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G101), .B1(new_n379), .B2(new_n380), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n350), .A3(KEYINPUT4), .ZN(new_n392));
  AND2_X1   g206(.A1(KEYINPUT0), .A2(G128), .ZN(new_n393));
  NOR2_X1   g207(.A1(KEYINPUT0), .A2(G128), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n364), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n364), .B2(new_n393), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(G101), .C1(new_n379), .C2(new_n380), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n343), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n334), .B1(new_n386), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n343), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n390), .B2(new_n399), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n382), .A2(new_n389), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n374), .A2(new_n387), .ZN(new_n407));
  AND4_X1   g221(.A1(new_n399), .A2(new_n406), .A3(new_n401), .A4(new_n407), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n405), .A2(new_n408), .A3(new_n333), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT82), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n350), .A2(new_n362), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n368), .A2(new_n355), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n404), .B(new_n372), .C1(new_n413), .C2(new_n374), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n384), .B1(new_n383), .B2(new_n343), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n402), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n333), .ZN(new_n417));
  INV_X1    g231(.A(new_n405), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n402), .A3(new_n334), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(G469), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n269), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n333), .B1(new_n405), .B2(new_n408), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n402), .B(new_n334), .C1(new_n414), .C2(new_n415), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n427), .B2(new_n423), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n330), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  OAI21_X1  g244(.A(G210), .B1(G237), .B2(G902), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n289), .A2(G119), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n289), .A2(KEYINPUT66), .A3(G119), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT66), .B1(new_n289), .B2(G119), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G113), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT2), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT2), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G113), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n444));
  INV_X1    g258(.A(G119), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(G116), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n289), .A2(KEYINPUT66), .A3(G119), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n433), .A3(new_n441), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n443), .A2(KEYINPUT67), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n448), .A2(new_n433), .A3(new_n441), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n441), .B1(new_n448), .B2(new_n433), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n392), .A2(new_n450), .A3(new_n454), .A4(new_n398), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n437), .B1(new_n456), .B2(new_n432), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n436), .B2(new_n456), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n382), .A2(new_n449), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n461), .A3(new_n459), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n396), .A2(G125), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n412), .B2(G125), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n467), .B(new_n469), .Z(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n467), .B(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n461), .B(KEYINPUT8), .Z(new_n477));
  INV_X1    g291(.A(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n457), .B1(new_n436), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n382), .A2(new_n449), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n458), .A2(new_n449), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n411), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(G902), .B1(new_n484), .B2(new_n464), .ZN(new_n485));
  AOI211_X1 g299(.A(KEYINPUT84), .B(new_n431), .C1(new_n473), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n473), .A2(new_n485), .ZN(new_n488));
  INV_X1    g302(.A(new_n431), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n473), .A2(new_n485), .A3(new_n431), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT84), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n429), .A2(new_n430), .A3(new_n487), .A4(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n328), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n309), .B1(G234), .B2(new_n269), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n445), .B2(G128), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n356), .A2(KEYINPUT23), .A3(G119), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n445), .A2(G128), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT73), .A4(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(G110), .A3(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT24), .B(G110), .Z(new_n505));
  XNOR2_X1  g319(.A(G119), .B(G128), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n244), .B2(new_n221), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n202), .A2(new_n195), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n500), .A2(G110), .B1(new_n505), .B2(new_n506), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n510), .A2(new_n221), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT77), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n252), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT77), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n221), .A3(new_n511), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(new_n517), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT77), .A3(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT25), .B1(new_n526), .B2(new_n269), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n528), .B(G902), .C1(new_n523), .C2(new_n525), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n495), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n495), .A2(G902), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n452), .A2(new_n453), .A3(new_n451), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT67), .B1(new_n443), .B2(new_n449), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n282), .A2(G137), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n337), .A2(G134), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n342), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n369), .A2(new_n541), .B1(new_n396), .B2(new_n343), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n454), .A2(KEYINPUT68), .A3(new_n450), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT69), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n537), .A2(new_n546), .A3(new_n542), .A4(new_n543), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n187), .A2(G210), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT27), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n369), .A2(KEYINPUT65), .A3(new_n541), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n396), .A2(new_n343), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT65), .B1(new_n369), .B2(new_n541), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n535), .A2(new_n536), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n542), .A2(KEYINPUT30), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n562));
  NAND4_X1  g376(.A1(new_n548), .A2(new_n552), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n561), .A2(new_n552), .A3(new_n545), .A4(new_n547), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n544), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n559), .B1(new_n556), .B2(new_n557), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n545), .A2(new_n547), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n569), .B2(KEYINPUT28), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n563), .B(new_n565), .C1(new_n570), .C2(new_n552), .ZN(new_n571));
  NOR2_X1   g385(.A1(G472), .A2(G902), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT32), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n572), .A2(KEYINPUT32), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n563), .A2(new_n565), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(KEYINPUT28), .ZN(new_n576));
  INV_X1    g390(.A(new_n567), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n552), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n574), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(KEYINPUT72), .A3(new_n574), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n573), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n537), .A2(new_n543), .ZN(new_n584));
  INV_X1    g398(.A(new_n542), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n545), .A2(new_n547), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n567), .B1(new_n587), .B2(KEYINPUT28), .ZN(new_n588));
  INV_X1    g402(.A(new_n552), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n548), .A2(new_n561), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n589), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n589), .B(new_n567), .C1(new_n569), .C2(KEYINPUT28), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT71), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n590), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n570), .A2(new_n552), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(KEYINPUT71), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n592), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n533), .B1(new_n583), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n494), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n273), .A2(new_n275), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n311), .A2(new_n312), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n314), .A3(new_n269), .ZN(new_n607));
  NAND2_X1  g421(.A1(G478), .A2(G902), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n606), .B(KEYINPUT33), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n314), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n490), .A2(new_n613), .A3(new_n491), .ZN(new_n614));
  INV_X1    g428(.A(new_n430), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n431), .B1(new_n473), .B2(new_n485), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(KEYINPUT96), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n612), .A2(new_n326), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n571), .A2(new_n269), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT94), .A3(G472), .ZN(new_n621));
  INV_X1    g435(.A(new_n533), .ZN(new_n622));
  NAND2_X1  g436(.A1(KEYINPUT94), .A2(G472), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n571), .A2(new_n269), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n621), .A2(new_n429), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT34), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  XNOR2_X1  g444(.A(new_n250), .B(new_n264), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n631), .A2(new_n271), .A3(new_n318), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n325), .A2(new_n632), .A3(new_n614), .A4(new_n617), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT98), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n638));
  INV_X1    g452(.A(new_n495), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n523), .A2(new_n525), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n528), .B1(new_n640), .B2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n526), .A2(KEYINPUT25), .A3(new_n269), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n524), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n531), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n638), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n530), .A2(KEYINPUT99), .A3(new_n646), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n621), .A2(new_n648), .A3(new_n624), .A4(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n328), .A2(new_n650), .A3(new_n493), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT37), .B(G110), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  NAND2_X1  g467(.A1(new_n648), .A2(new_n649), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n583), .B2(new_n601), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n320), .B1(new_n323), .B2(G900), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n632), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n429), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n618), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n656), .B(KEYINPUT39), .Z(new_n662));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n266), .A2(new_n274), .A3(new_n271), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n274), .B1(new_n266), .B2(new_n271), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n530), .A2(new_n646), .ZN(new_n668));
  NOR4_X1   g482(.A1(new_n667), .A2(new_n317), .A3(new_n615), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n593), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n589), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n269), .B1(new_n587), .B2(new_n552), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n583), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n492), .A2(new_n487), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n664), .A2(new_n669), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n583), .A2(new_n601), .ZN(new_n681));
  INV_X1    g495(.A(new_n654), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n659), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n611), .B(new_n656), .C1(new_n665), .C2(new_n666), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n684), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n655), .A3(KEYINPUT100), .A4(new_n659), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n423), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n427), .A2(new_n692), .ZN(new_n693));
  AOI211_X1 g507(.A(G902), .B(new_n691), .C1(new_n425), .C2(new_n426), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n330), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n602), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n619), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n633), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT102), .B(G116), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G18));
  NAND3_X1  g516(.A1(new_n695), .A2(new_n614), .A3(new_n617), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n328), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n655), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NAND3_X1  g520(.A1(new_n614), .A2(new_n318), .A3(new_n617), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT104), .B1(new_n667), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n707), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n605), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n572), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n587), .A2(KEYINPUT28), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n577), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n588), .A2(KEYINPUT103), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n589), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n563), .A2(new_n565), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n713), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(G472), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n571), .B2(new_n269), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n721), .A2(new_n533), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n325), .A3(new_n695), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n712), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT105), .B(G122), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G24));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n729));
  INV_X1    g543(.A(new_n668), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n721), .A2(new_n730), .A3(new_n723), .ZN(new_n731));
  INV_X1    g545(.A(new_n703), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n733), .B2(new_n684), .ZN(new_n734));
  INV_X1    g548(.A(new_n718), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n589), .B1(new_n588), .B2(KEYINPUT103), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n720), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n572), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n620), .A2(G472), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n668), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n703), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n734), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(new_n579), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(new_n573), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n598), .A2(KEYINPUT71), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n595), .A2(new_n596), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n590), .A4(new_n594), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n722), .B1(new_n749), .B2(new_n592), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n622), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(new_n622), .C1(new_n746), .C2(new_n750), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n417), .A2(new_n419), .A3(G469), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n330), .B1(new_n428), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n616), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n430), .B(new_n758), .C1(new_n760), .C2(new_n486), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n684), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n761), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n686), .A2(new_n602), .A3(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n755), .A2(new_n762), .B1(new_n764), .B2(new_n756), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n232), .ZN(G33));
  NAND4_X1  g580(.A1(new_n681), .A2(new_n763), .A3(new_n622), .A4(new_n657), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NOR2_X1   g582(.A1(new_n605), .A2(new_n610), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n605), .B2(new_n610), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n730), .B1(new_n621), .B2(new_n624), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT44), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(KEYINPUT44), .A3(new_n774), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n430), .B1(new_n760), .B2(new_n486), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n775), .B1(new_n780), .B2(KEYINPUT108), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT45), .B1(new_n410), .B2(new_n421), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(G469), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n424), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n791), .A2(new_n792), .B1(new_n423), .B2(new_n427), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n329), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n662), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n781), .A2(new_n798), .A3(new_n783), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n785), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  NOR4_X1   g615(.A1(new_n681), .A2(new_n684), .A3(new_n622), .A4(new_n777), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n329), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT47), .B1(new_n795), .B2(new_n329), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  AOI21_X1  g620(.A(new_n320), .B1(new_n770), .B2(new_n772), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n695), .A3(new_n778), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n754), .B2(new_n752), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT48), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(KEYINPUT48), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n807), .A2(new_n724), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(KEYINPUT119), .A3(new_n732), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT119), .B1(new_n812), .B2(new_n732), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n674), .A2(new_n533), .A3(new_n320), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n695), .A3(new_n778), .ZN(new_n817));
  OAI211_X1 g631(.A(G952), .B(new_n226), .C1(new_n817), .C2(new_n612), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n803), .A2(new_n804), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n693), .A2(new_n694), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n330), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n778), .A3(new_n812), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n808), .A2(new_n740), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n817), .A2(new_n605), .A3(new_n611), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n812), .A2(new_n615), .A3(new_n676), .A4(new_n695), .ZN(new_n829));
  XOR2_X1   g643(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n830));
  AND2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(KEYINPUT50), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n814), .B(new_n819), .C1(new_n828), .C2(new_n835), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT118), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT118), .B1(new_n831), .B2(new_n834), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n824), .A3(new_n827), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n740), .A2(new_n761), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n422), .A2(new_n428), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n271), .A2(new_n317), .A3(new_n656), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n329), .A3(new_n631), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n777), .A2(new_n846), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n686), .A2(new_n843), .B1(new_n655), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n842), .B1(new_n848), .B2(new_n767), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n610), .B1(new_n273), .B2(new_n275), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n763), .A2(new_n850), .A3(new_n656), .A4(new_n731), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n681), .A3(new_n682), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n842), .A2(new_n767), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n328), .A2(new_n650), .A3(new_n493), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n492), .A2(new_n487), .A3(new_n325), .A4(new_n430), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n625), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n667), .A3(new_n318), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n858), .A3(KEYINPUT110), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n273), .A2(new_n275), .A3(new_n318), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n861), .A2(new_n625), .A3(new_n856), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n651), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n602), .A2(new_n494), .B1(new_n857), .B2(new_n850), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n859), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n697), .A2(new_n700), .A3(new_n726), .A4(new_n705), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n765), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n730), .A2(new_n674), .A3(new_n656), .A4(new_n758), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n685), .A2(new_n687), .B1(new_n871), .B2(new_n712), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n734), .B2(new_n742), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n743), .A2(new_n660), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT112), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n743), .A2(new_n880), .A3(new_n660), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(KEYINPUT52), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n872), .A2(new_n874), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n866), .A2(new_n885), .A3(new_n887), .A4(new_n869), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n870), .A2(new_n884), .B1(new_n888), .B2(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n854), .B2(new_n865), .ZN(new_n893));
  INV_X1    g707(.A(new_n865), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n767), .A2(new_n851), .A3(new_n852), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT111), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n848), .A2(new_n842), .A3(new_n767), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n898), .A3(KEYINPUT114), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n868), .A2(new_n867), .A3(new_n765), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n743), .A2(new_n880), .A3(new_n660), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n880), .B1(new_n743), .B2(new_n660), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n904), .A2(new_n905), .B1(new_n875), .B2(new_n876), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n891), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n755), .A2(new_n762), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n764), .A2(new_n756), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n696), .A2(new_n619), .B1(new_n655), .B2(new_n704), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n633), .A2(new_n696), .B1(new_n712), .B2(new_n725), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(KEYINPUT53), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n894), .A2(new_n898), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n892), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n915), .A2(new_n884), .A3(KEYINPUT115), .A4(new_n899), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n888), .A2(new_n867), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n907), .A2(new_n916), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n841), .A2(new_n890), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(G952), .B2(G953), .ZN(new_n921));
  INV_X1    g735(.A(new_n674), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n622), .A2(new_n430), .A3(new_n329), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT49), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n821), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT49), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n676), .A2(new_n922), .A3(new_n769), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n226), .A2(G952), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT122), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n907), .A2(new_n916), .A3(new_n918), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n465), .A2(new_n472), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(new_n470), .Z(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n931), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n935), .A2(new_n939), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n935), .A2(KEYINPUT121), .A3(new_n939), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G51));
  INV_X1    g759(.A(new_n917), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n932), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(KEYINPUT123), .A3(new_n919), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n932), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n424), .B(KEYINPUT57), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n425), .A2(new_n426), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n932), .A2(G902), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n789), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n930), .B1(new_n955), .B2(new_n957), .ZN(G54));
  NAND2_X1  g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n956), .A2(new_n259), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n259), .B1(new_n956), .B2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n930), .ZN(G60));
  XOR2_X1   g777(.A(new_n608), .B(KEYINPUT59), .Z(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n890), .B2(new_n919), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n931), .B1(new_n965), .B2(new_n609), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n948), .A2(new_n950), .ZN(new_n967));
  INV_X1    g781(.A(new_n609), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n964), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n932), .A2(new_n645), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n932), .A2(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n931), .B(new_n973), .C1(new_n974), .C2(new_n526), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  NOR2_X1   g791(.A1(new_n868), .A2(new_n865), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n226), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  OAI21_X1  g796(.A(G953), .B1(new_n321), .B2(new_n468), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT127), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n936), .B1(G898), .B2(new_n226), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(new_n904), .A2(new_n688), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n797), .A2(new_n712), .A3(new_n755), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n805), .A3(new_n767), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n988), .A2(new_n990), .A3(new_n765), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n800), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n226), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n558), .A2(new_n560), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(new_n211), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(G900), .B2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n226), .B1(G227), .B2(G900), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n612), .A2(new_n861), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n602), .A3(new_n663), .A4(new_n778), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n805), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n904), .A2(new_n678), .A3(new_n688), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(KEYINPUT62), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n800), .B(new_n1005), .C1(KEYINPUT62), .C2(new_n1004), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1006), .A2(new_n226), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n998), .B(new_n1000), .C1(new_n1007), .C2(new_n995), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n995), .B1(new_n1006), .B2(new_n226), .ZN(new_n1009));
  INV_X1    g823(.A(new_n997), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1010), .B1(new_n992), .B2(new_n226), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n999), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1008), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n594), .A2(new_n564), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n889), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(G952), .B2(new_n226), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n670), .A2(new_n589), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n800), .A2(new_n991), .A3(new_n979), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(new_n1020), .B2(new_n1015), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1006), .B2(new_n980), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1018), .B(new_n1021), .C1(new_n1022), .C2(new_n671), .ZN(G57));
endmodule


