//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G244), .Z(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  AND3_X1   g0045(.A1(new_n245), .A2(KEYINPUT72), .A3(new_n213), .ZN(new_n246));
  AOI21_X1  g0046(.A(KEYINPUT72), .B1(new_n245), .B2(new_n213), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT24), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT85), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(new_n214), .A4(G87), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT78), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT78), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n260), .A3(G33), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n261), .A2(new_n214), .A3(G87), .A4(new_n251), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT85), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(new_n263), .A3(KEYINPUT22), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G87), .ZN(new_n267));
  OR4_X1    g0067(.A1(KEYINPUT22), .A2(new_n266), .A3(G20), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G107), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n250), .A2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G116), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n273), .A2(new_n274), .A3(new_n275), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n249), .B1(new_n269), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g0080(.A(KEYINPUT24), .B(new_n278), .C1(new_n264), .C2(new_n268), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n248), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n214), .A3(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n270), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT25), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n283), .A2(G1), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n288), .B(new_n290), .C1(new_n246), .C2(new_n247), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n286), .B1(G107), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n213), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  MUX2_X1   g0096(.A(G250), .B(G257), .S(G1698), .Z(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(new_n261), .A3(new_n251), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G294), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n289), .A2(G45), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT5), .A2(G41), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT5), .A2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(KEYINPUT69), .A2(G33), .A3(G41), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n294), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n308), .A3(G274), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G45), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G1), .ZN(new_n312));
  INV_X1    g0112(.A(new_n303), .ZN(new_n313));
  NOR2_X1   g0113(.A1(KEYINPUT5), .A2(G41), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n308), .A2(new_n315), .A3(G264), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n300), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G200), .B2(new_n317), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n282), .A2(new_n293), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  INV_X1    g0122(.A(new_n296), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n251), .A2(new_n265), .A3(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT70), .A3(G1698), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(G222), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n218), .B2(new_n328), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n323), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G41), .ZN(new_n335));
  AOI21_X1  g0135(.A(G1), .B1(new_n335), .B2(new_n311), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n213), .B1(new_n305), .B2(new_n295), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n307), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G226), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n289), .B1(G41), .B2(G45), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n340), .A2(new_n308), .A3(G274), .A4(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n322), .B1(new_n334), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n334), .A2(new_n322), .A3(new_n345), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT73), .B1(new_n248), .B2(new_n284), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT73), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n288), .C1(new_n246), .C2(new_n247), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n352), .A2(new_n354), .B1(new_n289), .B2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G50), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n203), .A2(G20), .ZN(new_n357));
  INV_X1    g0157(.A(G150), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G20), .A2(G33), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n276), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT8), .B(G58), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n357), .B1(new_n358), .B2(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n248), .B1(new_n202), .B2(new_n284), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n347), .A2(new_n366), .A3(new_n348), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n351), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT9), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n347), .A2(G200), .A3(new_n348), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT9), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT77), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n365), .A2(KEYINPUT77), .A3(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n349), .A2(G190), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n372), .A2(new_n373), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n370), .A3(new_n371), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT77), .B1(new_n365), .B2(new_n374), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n376), .B(KEYINPUT9), .C1(new_n356), .C2(new_n364), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT10), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n368), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G68), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n359), .A2(G50), .B1(G20), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G77), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n361), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n248), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT11), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n284), .A2(new_n388), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT12), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n246), .A2(new_n247), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n388), .B1(new_n289), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n288), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n248), .A2(new_n391), .A3(KEYINPUT11), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n394), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  MUX2_X1   g0201(.A(G226), .B(G232), .S(G1698), .Z(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n328), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n323), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n308), .A2(G238), .A3(new_n341), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n344), .A4(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n402), .A2(new_n328), .B1(G33), .B2(G97), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n344), .B(new_n408), .C1(new_n410), .C2(new_n296), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(G169), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n412), .A3(G179), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n413), .B2(G169), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n401), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n413), .A2(G200), .ZN(new_n420));
  INV_X1    g0220(.A(new_n401), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n318), .C2(new_n413), .ZN(new_n422));
  INV_X1    g0222(.A(new_n217), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n338), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n344), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n328), .A2(KEYINPUT74), .A3(G232), .A4(new_n331), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n328), .A2(G232), .A3(new_n331), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT74), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(G107), .B2(new_n266), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n327), .A2(new_n329), .ZN(new_n430));
  INV_X1    g0230(.A(G238), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n426), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n425), .B1(new_n432), .B2(new_n323), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n350), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n427), .A2(new_n428), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n266), .A2(G107), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n426), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n327), .B2(new_n329), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n323), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n425), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n366), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n390), .B1(new_n289), .B2(G20), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n397), .A2(new_n288), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n218), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n288), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G58), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT8), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT8), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G58), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT75), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n362), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n359), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT15), .B(G87), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(G20), .A2(new_n445), .B1(new_n458), .B2(new_n276), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n444), .B(new_n447), .C1(new_n460), .C2(new_n397), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n434), .A2(new_n442), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G200), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n439), .B2(new_n440), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT76), .B1(new_n464), .B2(new_n461), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n397), .B1(new_n456), .B2(new_n459), .ZN(new_n466));
  INV_X1    g0266(.A(new_n444), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n466), .A2(new_n467), .A3(new_n446), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT76), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n469), .C1(new_n433), .C2(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n433), .A2(G190), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n465), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n419), .A2(new_n422), .A3(new_n462), .A4(new_n472), .ZN(new_n473));
  MUX2_X1   g0273(.A(G223), .B(G226), .S(G1698), .Z(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n261), .A3(new_n251), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G87), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n296), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n479), .B(new_n296), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n338), .A2(G232), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n350), .A3(new_n344), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n344), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n366), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT81), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(G58), .A2(G68), .ZN(new_n488));
  OAI21_X1  g0288(.A(G20), .B1(new_n488), .B2(new_n201), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n359), .A2(G159), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(KEYINPUT79), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT79), .B1(new_n489), .B2(new_n490), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n261), .A2(new_n251), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT7), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n214), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G68), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n495), .B2(new_n214), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT16), .B(new_n494), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT16), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n496), .A2(G20), .ZN(new_n502));
  AOI21_X1  g0302(.A(G33), .B1(new_n258), .B2(new_n260), .ZN(new_n503));
  INV_X1    g0303(.A(new_n265), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n496), .B1(new_n328), .B2(G20), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n388), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n489), .A2(new_n490), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT79), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n491), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n501), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n500), .A2(new_n248), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n288), .A2(new_n362), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n355), .B2(new_n362), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n475), .A2(new_n476), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n323), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n479), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n517), .B(new_n485), .C1(new_n522), .C2(new_n482), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n487), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT18), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT18), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n487), .A2(new_n516), .A3(new_n523), .A4(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n463), .B1(new_n484), .B2(new_n477), .ZN(new_n528));
  INV_X1    g0328(.A(new_n484), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n318), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(new_n513), .A3(new_n515), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT82), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n513), .A3(new_n515), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n525), .A2(new_n527), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n387), .A2(new_n473), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G238), .A2(G1698), .ZN(new_n541));
  INV_X1    g0341(.A(G244), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(G1698), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n261), .A3(new_n251), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n296), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n301), .A2(KEYINPUT83), .ZN(new_n547));
  OR3_X1    g0347(.A1(new_n311), .A2(KEYINPUT83), .A3(G1), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n308), .A2(G250), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n308), .A2(G274), .A3(new_n312), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G190), .ZN(new_n553));
  OAI21_X1  g0353(.A(G200), .B1(new_n546), .B2(new_n551), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n276), .A2(new_n555), .A3(G97), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n267), .B1(new_n404), .B2(new_n214), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n558), .B2(new_n555), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n261), .A2(new_n214), .A3(G68), .A4(new_n251), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n248), .B1(new_n284), .B2(new_n457), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n292), .A2(G87), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n553), .A2(new_n554), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n292), .A2(new_n458), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n552), .A2(new_n350), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n366), .B1(new_n546), .B2(new_n551), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n542), .A2(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n495), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(KEYINPUT4), .A2(G244), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n251), .A2(new_n265), .A3(new_n575), .A4(new_n331), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n251), .A2(new_n265), .A3(G250), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G283), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n296), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n308), .A2(new_n315), .A3(G257), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n309), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n350), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n366), .B1(new_n580), .B2(new_n582), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n270), .B1(new_n505), .B2(new_n506), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT6), .ZN(new_n587));
  INV_X1    g0387(.A(G97), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n587), .A2(new_n588), .A3(G107), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n591), .A2(new_n214), .B1(new_n390), .B2(new_n360), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n248), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n288), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n292), .B2(G97), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n584), .A2(new_n585), .A3(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n580), .A2(G190), .A3(new_n582), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT4), .B1(new_n254), .B2(new_n572), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n323), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n582), .ZN(new_n602));
  AOI21_X1  g0402(.A(G200), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n593), .B(new_n595), .C1(new_n598), .C2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n570), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n292), .A2(G116), .ZN(new_n606));
  INV_X1    g0406(.A(new_n287), .ZN(new_n607));
  INV_X1    g0407(.A(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G20), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n578), .B(new_n214), .C1(G33), .C2(new_n588), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n245), .A2(new_n213), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n609), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT20), .A4(new_n609), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  MUX2_X1   g0419(.A(G257), .B(G264), .S(G1698), .Z(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n261), .A3(new_n251), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n266), .A2(G303), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n296), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n308), .A2(new_n315), .A3(G270), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT84), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n309), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n309), .B2(new_n625), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n624), .B(G190), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n309), .A2(new_n625), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT84), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n309), .A2(new_n625), .A3(new_n626), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n623), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n619), .B(new_n629), .C1(new_n633), .C2(new_n463), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n623), .A2(new_n350), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n618), .B(new_n635), .C1(new_n627), .C2(new_n628), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n366), .B1(new_n606), .B2(new_n617), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT21), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n637), .B2(new_n638), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n634), .B(new_n636), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n282), .A2(new_n293), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n317), .A2(G169), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n317), .A2(new_n350), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n642), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n321), .A2(new_n540), .A3(new_n605), .A4(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n569), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n584), .A2(new_n596), .A3(new_n585), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n570), .A2(new_n651), .A3(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n564), .A2(new_n569), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n597), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n650), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n604), .A2(new_n597), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n321), .A2(new_n657), .A3(new_n570), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n643), .B2(new_n647), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n540), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n525), .A2(new_n527), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n462), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n422), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n419), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n535), .A2(new_n537), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n381), .A2(new_n386), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n368), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n671), .ZN(G369));
  INV_X1    g0472(.A(new_n642), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n607), .A2(KEYINPUT27), .A3(G20), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT27), .B1(new_n607), .B2(G20), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n673), .B1(new_n619), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n659), .A2(new_n618), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT87), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT87), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(new_n684), .A3(new_n681), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(KEYINPUT88), .B(G330), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n646), .B1(new_n282), .B2(new_n293), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n643), .A2(new_n678), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n321), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n679), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n659), .A2(new_n679), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n693), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n207), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n557), .A2(new_n267), .A3(new_n608), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n702), .A2(new_n703), .A3(new_n289), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n212), .B2(new_n702), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  NAND2_X1  g0506(.A1(new_n661), .A2(new_n679), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n605), .B(new_n321), .C1(new_n689), .C2(new_n659), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n678), .B1(new_n709), .B2(new_n656), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n648), .A2(new_n321), .A3(new_n605), .A4(new_n679), .ZN(new_n714));
  NOR4_X1   g0514(.A1(new_n583), .A2(new_n317), .A3(G179), .A4(new_n552), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n638), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n601), .B(new_n602), .C1(new_n627), .C2(new_n628), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n300), .A2(new_n316), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n552), .A2(new_n718), .A3(new_n635), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT89), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT30), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  OAI211_X1 g0522(.A(KEYINPUT89), .B(new_n722), .C1(new_n717), .C2(new_n719), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n716), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n678), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n714), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n687), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n713), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n706), .B1(new_n732), .B2(G1), .ZN(G364));
  OR2_X1    g0533(.A1(new_n686), .A2(new_n687), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n283), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n289), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n702), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n734), .A2(new_n688), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n701), .A2(new_n266), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G355), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G116), .B2(new_n207), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n701), .B(new_n254), .C1(new_n311), .C2(new_n212), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n243), .A2(G45), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OR3_X1    g0546(.A1(KEYINPUT90), .A2(G13), .A3(G33), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT90), .B1(G13), .B2(G33), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n213), .B1(G20), .B2(new_n366), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n738), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n214), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n267), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n214), .A2(new_n350), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n756), .A2(new_n318), .A3(G200), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n388), .B1(new_n763), .B2(new_n270), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n760), .A2(new_n318), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n758), .B(new_n764), .C1(G50), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n756), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G159), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT32), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n318), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n214), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n770), .A2(KEYINPUT32), .B1(new_n774), .B2(G97), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n759), .A2(G190), .A3(new_n463), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n328), .B1(new_n776), .B2(new_n448), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n759), .A2(new_n767), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(new_n445), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n766), .A2(new_n771), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n765), .B(KEYINPUT91), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n757), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n774), .A2(G294), .B1(new_n785), .B2(G303), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  INV_X1    g0587(.A(new_n763), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n761), .A2(new_n787), .B1(new_n788), .B2(G283), .ZN(new_n789));
  INV_X1    g0589(.A(new_n776), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G322), .B1(new_n779), .B2(G311), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n328), .B1(new_n769), .B2(G329), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n786), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n781), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT92), .ZN(new_n795));
  INV_X1    g0595(.A(new_n752), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n794), .B2(KEYINPUT92), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n755), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n751), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n682), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT93), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n740), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NOR2_X1   g0603(.A1(new_n462), .A2(new_n678), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n461), .A2(new_n678), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n472), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(new_n806), .B2(new_n462), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n707), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n661), .A2(new_n679), .A3(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n738), .B1(new_n811), .B2(new_n730), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n730), .B2(new_n811), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n750), .A2(new_n796), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n738), .B1(new_n814), .B2(G77), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  INV_X1    g0616(.A(new_n765), .ZN(new_n817));
  INV_X1    g0617(.A(G303), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n816), .A2(new_n762), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G107), .B2(new_n785), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n776), .A2(new_n821), .B1(new_n768), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n328), .B(new_n823), .C1(G116), .C2(new_n779), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n763), .A2(new_n267), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G97), .B2(new_n774), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n820), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n790), .A2(G143), .B1(new_n779), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n817), .B2(new_n829), .C1(new_n358), .C2(new_n762), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  AOI21_X1  g0631(.A(new_n495), .B1(G132), .B2(new_n769), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n832), .A2(KEYINPUT94), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n763), .A2(new_n388), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n773), .A2(new_n448), .B1(new_n757), .B2(new_n202), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(KEYINPUT94), .B2(new_n832), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n827), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n815), .B1(new_n838), .B2(new_n752), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT95), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n750), .B2(new_n807), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n813), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  INV_X1    g0643(.A(new_n591), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT35), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(KEYINPUT35), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(G116), .A3(new_n215), .A4(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT36), .Z(new_n848));
  OR3_X1    g0648(.A1(new_n211), .A2(new_n218), .A3(new_n488), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n202), .A2(G68), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n289), .B(G13), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT99), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n419), .A2(new_n678), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n500), .A2(new_n248), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT7), .B1(new_n254), .B2(G20), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(G68), .A3(new_n497), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT16), .B1(new_n858), .B2(new_n494), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n515), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n676), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n538), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n487), .A3(new_n523), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n532), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n516), .A2(new_n861), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n524), .A2(new_n868), .A3(new_n532), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n864), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n869), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n538), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n524), .A2(new_n532), .A3(new_n869), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n870), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT97), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n538), .A2(new_n875), .B1(new_n878), .B2(new_n870), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT97), .B1(new_n884), .B2(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n874), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n864), .B2(new_n871), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n873), .B1(new_n888), .B2(new_n872), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT98), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n538), .A2(new_n863), .B1(new_n867), .B2(new_n870), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT39), .B1(new_n892), .B2(KEYINPUT38), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n894));
  AOI211_X1 g0694(.A(KEYINPUT97), .B(KEYINPUT38), .C1(new_n876), .C2(new_n879), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n872), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT39), .B1(new_n897), .B2(new_n887), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT98), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n855), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n804), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n810), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT96), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n401), .A2(new_n678), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n419), .A2(new_n422), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n419), .B2(new_n422), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT96), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n810), .A2(new_n908), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n897), .A2(new_n887), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n910), .A2(new_n911), .B1(new_n664), .B2(new_n861), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n853), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n890), .B1(new_n886), .B2(new_n889), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n896), .A2(KEYINPUT98), .A3(new_n898), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n854), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n917), .A2(KEYINPUT99), .A3(new_n912), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n540), .B1(new_n708), .B2(new_n712), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n671), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n807), .B1(new_n905), .B2(new_n906), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n729), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n923), .B1(new_n911), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(KEYINPUT100), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT100), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n929), .A3(new_n729), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(KEYINPUT40), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n897), .B1(new_n885), .B2(new_n883), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n540), .A2(new_n729), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n687), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n922), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n289), .B2(new_n735), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n922), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n852), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NOR2_X1   g0741(.A1(new_n694), .A2(new_n697), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n596), .A2(new_n678), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n657), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n651), .A2(new_n678), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n689), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n597), .B1(new_n948), .B2(new_n944), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n947), .A2(KEYINPUT42), .B1(new_n679), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT42), .B2(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n562), .A2(new_n563), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n678), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n570), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT101), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT101), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(new_n569), .C2(new_n953), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT102), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n951), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n960), .B1(new_n951), .B2(new_n961), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n695), .A2(new_n946), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n702), .B(KEYINPUT41), .Z(new_n967));
  INV_X1    g0767(.A(new_n946), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n698), .A2(KEYINPUT103), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT103), .B1(new_n698), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n698), .A2(new_n968), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT44), .Z(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(new_n695), .ZN(new_n978));
  INV_X1    g0778(.A(new_n942), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n694), .A2(new_n697), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n688), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n688), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n731), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n977), .A2(new_n695), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n967), .B1(new_n986), .B2(new_n732), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n965), .B(new_n966), .C1(new_n987), .C2(new_n737), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n753), .B1(new_n207), .B2(new_n457), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n254), .A2(new_n701), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n989), .B1(new_n235), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n782), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(G143), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n778), .A2(new_n202), .B1(new_n768), .B2(new_n829), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n266), .B(new_n994), .C1(G150), .C2(new_n790), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n774), .A2(G68), .B1(new_n788), .B2(new_n445), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n761), .A2(G159), .B1(new_n785), .B2(G58), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT107), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n757), .A2(new_n608), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n762), .A2(new_n821), .B1(KEYINPUT46), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT46), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT105), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n763), .A2(new_n588), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT106), .B(G317), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n495), .B1(new_n768), .B2(new_n1005), .C1(new_n818), .C2(new_n776), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(new_n992), .C2(G311), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1002), .A2(KEYINPUT105), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n773), .A2(new_n270), .B1(new_n778), .B2(new_n816), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT104), .Z(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n999), .B1(new_n1003), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n739), .B(new_n991), .C1(new_n1013), .C2(new_n752), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n799), .B2(new_n957), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n988), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n694), .A2(new_n751), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n741), .A2(new_n703), .B1(new_n270), .B2(new_n701), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n453), .A2(new_n455), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(G50), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT50), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n311), .B1(new_n388), .B2(new_n390), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n703), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n232), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n990), .B1(new_n1024), .B2(new_n311), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1018), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n739), .B1(new_n1026), .B2(new_n753), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n757), .A2(new_n218), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n452), .B2(new_n761), .ZN(new_n1029));
  INV_X1    g0829(.A(G159), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n817), .C1(new_n457), .C2(new_n773), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n790), .A2(G50), .B1(new_n779), .B2(G68), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n358), .B2(new_n768), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1031), .A2(new_n495), .A3(new_n1004), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1005), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n790), .A2(new_n1035), .B1(new_n779), .B2(G303), .ZN(new_n1036));
  INV_X1    g0836(.A(G322), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1036), .B1(new_n822), .B2(new_n762), .C1(new_n782), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n774), .A2(G283), .B1(new_n785), .B2(G294), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n495), .B1(new_n608), .B2(new_n763), .C1(new_n783), .C2(new_n768), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1044), .B2(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1034), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1017), .B(new_n1027), .C1(new_n796), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n983), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT108), .B1(new_n1050), .B2(new_n737), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1050), .A2(KEYINPUT108), .A3(new_n737), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n983), .A2(new_n731), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT109), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n984), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n702), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1053), .A2(KEYINPUT109), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .C1(new_n1056), .C2(new_n1057), .ZN(G393));
  NAND3_X1  g0858(.A1(new_n978), .A2(new_n737), .A3(new_n985), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n240), .A2(new_n990), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n753), .C1(new_n588), .C2(new_n207), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT110), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT110), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n738), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n817), .A2(new_n358), .B1(new_n1030), .B2(new_n776), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n785), .A2(G68), .B1(new_n769), .B2(G143), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT111), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT111), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n495), .B(new_n825), .C1(G77), .C2(new_n774), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1019), .A2(new_n778), .B1(new_n762), .B2(new_n202), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT112), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G317), .A2(new_n765), .B1(new_n790), .B2(G311), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n762), .A2(new_n818), .B1(new_n763), .B2(new_n270), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n266), .B1(new_n768), .B2(new_n1037), .C1(new_n821), .C2(new_n778), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n773), .A2(new_n608), .B1(new_n757), .B2(new_n816), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1071), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1064), .B1(new_n752), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n799), .B2(new_n946), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n986), .A2(new_n702), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n984), .B1(new_n978), .B2(new_n985), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1059), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(G390));
  NAND2_X1  g0885(.A1(new_n910), .A2(new_n854), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n915), .A3(new_n916), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n932), .A2(new_n855), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n905), .A2(new_n906), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n804), .B1(new_n710), .B2(new_n807), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT113), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n729), .A2(G330), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n924), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n925), .A2(new_n729), .A3(KEYINPUT113), .A4(G330), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n729), .A2(new_n907), .A3(new_n687), .A4(new_n807), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1087), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n736), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n738), .B1(new_n814), .B2(new_n452), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n891), .A2(new_n899), .A3(new_n750), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n270), .A2(new_n762), .B1(new_n817), .B2(new_n816), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n266), .B1(new_n768), .B2(new_n821), .C1(new_n588), .C2(new_n778), .ZN(new_n1106));
  OR4_X1    g0906(.A1(new_n758), .A2(new_n1105), .A3(new_n834), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n773), .A2(new_n390), .B1(new_n776), .B2(new_n608), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT118), .Z(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n761), .A2(G137), .B1(new_n779), .B2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT117), .Z(new_n1113));
  INV_X1    g0913(.A(G125), .ZN(new_n1114));
  INV_X1    g0914(.A(G132), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n328), .B1(new_n768), .B2(new_n1114), .C1(new_n776), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n785), .A2(G150), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(KEYINPUT53), .B2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n773), .A2(new_n1030), .B1(new_n763), .B2(new_n202), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G128), .B2(new_n765), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(KEYINPUT53), .C2(new_n1117), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1107), .A2(new_n1109), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1103), .B(new_n1104), .C1(new_n752), .C2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1102), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n729), .A2(new_n687), .A3(new_n807), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1089), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1095), .A2(new_n1096), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n909), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n908), .B1(new_n810), .B2(new_n901), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT114), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n729), .A2(G330), .A3(new_n807), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n907), .ZN(new_n1135));
  OAI211_X1 g0935(.A(KEYINPUT114), .B(new_n1089), .C1(new_n1094), .C2(new_n808), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1099), .A2(new_n1090), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n540), .A2(G330), .A3(new_n729), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n920), .A2(new_n1140), .A3(new_n671), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT115), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1144), .B(new_n1141), .C1(new_n1132), .C2(new_n1138), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1125), .B(new_n702), .C1(new_n1101), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1101), .A2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1098), .B(new_n1100), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1125), .B1(new_n1150), .B2(new_n702), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1124), .B1(new_n1149), .B2(new_n1151), .ZN(G378));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1087), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1087), .A2(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1144), .B1(new_n1157), .B2(new_n1141), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1139), .A2(KEYINPUT115), .A3(new_n1142), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1141), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n927), .B(G330), .C1(new_n931), .C2(new_n932), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n369), .A2(new_n676), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n387), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n387), .A2(new_n1164), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1167), .B(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1162), .B(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n914), .B2(new_n918), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n900), .A2(new_n853), .A3(new_n913), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT99), .B1(new_n917), .B2(new_n912), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1162), .A2(new_n1170), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1162), .A2(new_n1170), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1153), .B1(new_n1161), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1142), .B1(new_n1101), .B2(new_n1146), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1177), .A4(new_n1172), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n702), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1172), .A2(new_n1177), .A3(new_n737), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1170), .A2(new_n749), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n738), .B1(new_n814), .B2(G50), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1114), .A2(new_n817), .B1(new_n762), .B2(new_n1115), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n790), .A2(G128), .B1(new_n779), .B2(G137), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n757), .B2(new_n1110), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G150), .C2(new_n774), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n788), .A2(G159), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n790), .A2(G107), .B1(new_n769), .B2(G283), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n457), .B2(new_n778), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1028), .B(new_n1197), .C1(G68), .C2(new_n774), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n817), .A2(new_n608), .B1(new_n763), .B2(new_n448), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G97), .B2(new_n761), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1198), .A2(new_n335), .A3(new_n495), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G50), .B1(new_n250), .B2(new_n335), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n254), .B2(G41), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1195), .A2(new_n1203), .A3(new_n1204), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1185), .B1(new_n1207), .B2(new_n752), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1184), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1183), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1182), .A2(new_n1211), .ZN(G375));
  OAI21_X1  g1012(.A(new_n738), .B1(new_n814), .B2(G68), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n817), .A2(new_n821), .B1(new_n763), .B2(new_n390), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G97), .B2(new_n785), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n776), .A2(new_n816), .B1(new_n768), .B2(new_n818), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n328), .B(new_n1216), .C1(G107), .C2(new_n779), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n458), .A2(new_n774), .B1(new_n761), .B2(G116), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n778), .A2(new_n358), .B1(new_n768), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G137), .B2(new_n790), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G50), .A2(new_n774), .B1(new_n761), .B2(new_n1111), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n765), .A2(G132), .B1(new_n785), .B2(G159), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n495), .B1(G58), .B2(new_n788), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1213), .B1(new_n1227), .B2(new_n752), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n907), .B2(new_n750), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1157), .A2(new_n736), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT120), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1231), .B2(new_n1230), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1157), .A2(new_n1141), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n967), .B(KEYINPUT119), .Z(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1146), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(G381));
  NOR4_X1   g1038(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1239));
  INV_X1    g1039(.A(G390), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G387), .A2(new_n1241), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1042(.A1(new_n677), .A2(G213), .ZN(new_n1243));
  OR2_X1    g1043(.A1(G378), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G375), .C2(new_n1244), .ZN(G409));
  NAND3_X1  g1045(.A1(new_n988), .A2(new_n1015), .A3(G390), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT124), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n988), .A2(new_n1248), .A3(new_n1015), .A4(G390), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(new_n1240), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(G393), .B(new_n802), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1253), .B(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1250), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1246), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1256), .A2(new_n1252), .A3(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1160), .A2(new_n1234), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n702), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT122), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1234), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1263), .B2(KEYINPUT60), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1260), .B(new_n1264), .C1(KEYINPUT60), .C2(new_n1263), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(G384), .A3(new_n1233), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G384), .B1(new_n1265), .B2(new_n1233), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1182), .A2(G378), .A3(new_n1211), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1180), .A2(new_n1177), .A3(new_n1172), .A4(new_n1236), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT121), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1210), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1178), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1274), .A2(KEYINPUT121), .A3(new_n1180), .A4(new_n1236), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G378), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1243), .B(new_n1269), .C1(new_n1270), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT123), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1211), .A3(new_n1275), .ZN(new_n1280));
  INV_X1    g1080(.A(G378), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1182), .A2(G378), .A3(new_n1211), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1243), .A4(new_n1269), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1278), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1243), .B1(new_n1270), .B2(new_n1276), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT126), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT126), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(new_n1292), .A3(new_n1243), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1293), .A3(KEYINPUT63), .A4(new_n1269), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1295));
  XOR2_X1   g1095(.A(new_n1269), .B(new_n1295), .Z(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1290), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1259), .A2(new_n1289), .A3(new_n1294), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1296), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1269), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1291), .A2(new_n1293), .A3(new_n1305), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(KEYINPUT127), .A2(new_n1306), .B1(new_n1287), .B2(new_n1304), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n1306), .A2(KEYINPUT127), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1302), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1298), .B1(new_n1309), .B2(new_n1259), .ZN(G405));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1281), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1283), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1303), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1259), .B(new_n1313), .ZN(G402));
endmodule


