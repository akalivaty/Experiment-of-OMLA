//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G101), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(KEYINPUT78), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n190), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G107), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(KEYINPUT76), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n191), .A2(KEYINPUT76), .A3(KEYINPUT3), .A4(G104), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n204), .A2(KEYINPUT84), .ZN(new_n205));
  INV_X1    g019(.A(G113), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT5), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT5), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT2), .B(G113), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n211), .A2(new_n213), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n216), .ZN(new_n218));
  XNOR2_X1  g032(.A(G110), .B(G122), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT8), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  OR2_X1    g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G143), .B(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G125), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n222), .A2(G143), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n226), .A2(new_n234), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n223), .A2(new_n225), .A3(new_n237), .A4(G128), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n233), .B1(G125), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G224), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT7), .B1(new_n241), .B2(G953), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n240), .A2(new_n243), .A3(new_n242), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n240), .B2(new_n242), .ZN(new_n245));
  OAI221_X1 g059(.A(new_n221), .B1(new_n240), .B2(new_n242), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n194), .B1(new_n200), .B2(new_n202), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n215), .A2(new_n212), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n207), .A2(G116), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n214), .B1(new_n209), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n191), .A2(KEYINPUT76), .A3(G104), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n201), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n190), .B1(new_n259), .B2(new_n194), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n255), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n247), .A2(G101), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n197), .B1(new_n258), .B2(new_n201), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(new_n248), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT77), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n254), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n196), .A2(new_n203), .A3(new_n216), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n219), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n189), .B1(new_n246), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n274));
  INV_X1    g088(.A(new_n219), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n249), .A2(new_n253), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n261), .B1(new_n255), .B2(new_n260), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n263), .A2(KEYINPUT77), .A3(new_n265), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n274), .B(new_n275), .C1(new_n279), .C2(new_n268), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n267), .A2(new_n269), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n274), .B1(new_n282), .B2(new_n275), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT82), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n278), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n268), .B1(new_n285), .B2(new_n254), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT81), .B1(new_n286), .B2(new_n219), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n286), .B2(new_n219), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .A4(new_n280), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n286), .A2(new_n219), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n241), .A2(G953), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n240), .B(new_n295), .ZN(new_n296));
  AND4_X1   g110(.A1(KEYINPUT83), .A2(new_n292), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n294), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n284), .B2(new_n291), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT83), .B1(new_n299), .B2(new_n296), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n273), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n302), .B(new_n273), .C1(new_n297), .C2(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n188), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT20), .ZN(new_n307));
  NOR2_X1   g121(.A1(G475), .A2(G902), .ZN(new_n308));
  XNOR2_X1  g122(.A(G113), .B(G122), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT87), .B(G104), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n222), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n316), .A2(KEYINPUT73), .A3(G125), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n312), .B2(KEYINPUT73), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n222), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G237), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G214), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n224), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT18), .A2(G131), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(G131), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n333), .A3(new_n326), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(KEYINPUT88), .A3(new_n332), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n312), .A2(KEYINPUT73), .ZN(new_n340));
  INV_X1    g154(.A(new_n317), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(KEYINPUT16), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G146), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n222), .A3(new_n345), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n327), .A2(KEYINPUT17), .A3(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n311), .B(new_n330), .C1(new_n339), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n346), .A2(G146), .B1(new_n331), .B2(new_n334), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n318), .A2(KEYINPUT86), .A3(KEYINPUT19), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT19), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n313), .A2(new_n314), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT86), .B1(new_n318), .B2(KEYINPUT19), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(G146), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n311), .B1(new_n359), .B2(new_n330), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n307), .B(new_n308), .C1(new_n352), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n308), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT89), .B1(new_n352), .B2(new_n360), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n357), .ZN(new_n365));
  INV_X1    g179(.A(new_n354), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n222), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n368), .A2(new_n353), .B1(new_n320), .B2(new_n329), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n364), .B(new_n351), .C1(new_n369), .C2(new_n311), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n362), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n361), .B1(new_n371), .B2(new_n307), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n330), .B1(new_n339), .B2(new_n350), .ZN(new_n373));
  INV_X1    g187(.A(new_n311), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n351), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n189), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(G475), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G478), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT15), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n383));
  INV_X1    g197(.A(G116), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(G122), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT90), .A3(G116), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n385), .A2(new_n387), .B1(new_n384), .B2(G122), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(KEYINPUT14), .B2(new_n191), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n224), .B2(G128), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n234), .A2(KEYINPUT92), .A3(G143), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n224), .A2(G128), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n388), .A2(new_n191), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n385), .B2(new_n387), .ZN(new_n401));
  OAI221_X1 g215(.A(new_n389), .B1(new_n397), .B2(new_n398), .C1(new_n399), .C2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n388), .B(new_n191), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT13), .B1(new_n224), .B2(G128), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT93), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(new_n224), .A3(KEYINPUT13), .A4(G128), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n393), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G134), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n403), .A2(new_n412), .A3(new_n396), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(G217), .A3(new_n322), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n402), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT94), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI211_X1 g237(.A(KEYINPUT94), .B(G902), .C1(new_n418), .C2(new_n420), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n382), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n402), .A2(new_n413), .A3(new_n419), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n419), .B1(new_n402), .B2(new_n413), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT94), .B1(new_n428), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n382), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G952), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  NAND2_X1  g248(.A1(G234), .A2(G237), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(G902), .A3(G953), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G898), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n380), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  INV_X1    g257(.A(new_n232), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n249), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n277), .B2(new_n278), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT11), .B1(new_n448), .B2(G134), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT64), .B(G137), .ZN(new_n452));
  AND2_X1   g266(.A1(KEYINPUT11), .A2(G134), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT65), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n448), .A2(KEYINPUT64), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G137), .ZN(new_n457));
  AND4_X1   g271(.A1(KEYINPUT65), .A2(new_n455), .A3(new_n457), .A4(new_n453), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n451), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n457), .A3(new_n453), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n452), .A2(KEYINPUT65), .A3(new_n453), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n333), .A3(new_n451), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n204), .ZN(new_n469));
  INV_X1    g283(.A(new_n239), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n238), .A2(KEYINPUT79), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT79), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n230), .A2(new_n474), .A3(new_n237), .A4(G128), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n236), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n196), .A2(new_n476), .A3(new_n203), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n469), .A2(new_n472), .B1(new_n477), .B2(new_n471), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n447), .A2(new_n468), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT78), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n195), .B(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n470), .B1(new_n481), .B2(new_n264), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n482), .A2(KEYINPUT80), .A3(new_n477), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n204), .A2(new_n484), .A3(new_n470), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n467), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT12), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(KEYINPUT80), .A3(new_n477), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n467), .A4(new_n485), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G140), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n322), .A2(G227), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AND4_X1   g308(.A1(new_n479), .A2(new_n487), .A3(new_n490), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n469), .A2(new_n472), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n477), .A2(new_n471), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n467), .B1(new_n498), .B2(new_n446), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n494), .B1(new_n499), .B2(new_n479), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n443), .B(new_n189), .C1(new_n495), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(G469), .A2(G902), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n479), .A2(new_n487), .A3(new_n490), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n493), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n479), .A3(new_n494), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(G469), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n207), .B2(G128), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n234), .A2(KEYINPUT23), .A3(G119), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n510), .C1(G119), .C2(new_n234), .ZN(new_n511));
  XNOR2_X1  g325(.A(G119), .B(G128), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT24), .B(G110), .Z(new_n513));
  OAI22_X1  g327(.A1(new_n511), .A2(G110), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n347), .A2(new_n315), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n347), .A2(new_n348), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(G110), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n512), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n515), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT75), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G137), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n515), .B(new_n525), .C1(new_n516), .C2(new_n520), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G234), .ZN(new_n532));
  OAI21_X1  g346(.A(G217), .B1(new_n532), .B2(G902), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT71), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n529), .B2(new_n530), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n527), .A2(new_n528), .ZN(new_n536));
  INV_X1    g350(.A(new_n534), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G902), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n531), .A2(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n507), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n232), .B1(new_n460), .B2(new_n466), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n449), .A2(new_n450), .ZN(new_n544));
  AOI211_X1 g358(.A(G131), .B(new_n544), .C1(new_n463), .C2(new_n464), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n450), .B1(new_n452), .B2(G134), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G131), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n239), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n253), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n333), .B1(new_n465), .B2(new_n451), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n444), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n250), .A2(new_n252), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n466), .A2(new_n239), .A3(new_n547), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n555), .A3(KEYINPUT69), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n557), .B(new_n253), .C1(new_n543), .C2(new_n549), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(KEYINPUT28), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n543), .B2(new_n549), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(KEYINPUT68), .A3(new_n554), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n553), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n325), .A2(G210), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n566), .B(KEYINPUT27), .Z(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT26), .B(G101), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND4_X1  g383(.A1(new_n559), .A2(new_n565), .A3(KEYINPUT29), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT70), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT66), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n545), .B2(new_n548), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n466), .A2(KEYINPUT66), .A3(new_n239), .A4(new_n547), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n552), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(new_n253), .ZN(new_n576));
  INV_X1    g390(.A(new_n555), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT28), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n569), .A3(new_n565), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n554), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n253), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n555), .ZN(new_n584));
  INV_X1    g398(.A(new_n569), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT29), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n189), .ZN(new_n589));
  OAI21_X1  g403(.A(G472), .B1(new_n571), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G472), .A2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n569), .B1(new_n578), .B2(new_n565), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT31), .ZN(new_n594));
  AND4_X1   g408(.A1(new_n594), .A2(new_n583), .A3(new_n555), .A4(new_n569), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n583), .A2(new_n555), .A3(new_n569), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT67), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n583), .A2(KEYINPUT67), .A3(new_n555), .A4(new_n569), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT31), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n592), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT32), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(KEYINPUT32), .B(new_n592), .C1(new_n596), .C2(new_n601), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n590), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n306), .A2(new_n442), .A3(new_n542), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  INV_X1    g422(.A(new_n441), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n428), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n426), .B2(new_n427), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(G478), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n421), .A2(new_n381), .ZN(new_n614));
  NAND2_X1  g428(.A1(G478), .A2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT95), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT95), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n613), .A2(new_n618), .A3(new_n614), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n380), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n306), .A2(new_n609), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n596), .A2(new_n601), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n189), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n627), .A2(new_n541), .A3(new_n602), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n306), .A2(new_n629), .A3(new_n609), .A4(new_n622), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n624), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n363), .A2(new_n370), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n308), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT20), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n371), .A2(new_n307), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n378), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n432), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n306), .A2(new_n609), .A3(new_n628), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR2_X1   g458(.A1(new_n627), .A2(new_n602), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n507), .A2(new_n540), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n531), .A2(new_n535), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n521), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n538), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n306), .A2(new_n442), .A3(new_n645), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT98), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND3_X1  g470(.A1(new_n606), .A2(new_n646), .A3(new_n651), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT99), .B(G900), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n439), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n436), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n639), .A2(new_n432), .A3(new_n661), .ZN(new_n662));
  AOI211_X1 g476(.A(new_n188), .B(new_n662), .C1(new_n304), .C2(new_n305), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  NAND2_X1  g479(.A1(new_n304), .A2(new_n305), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT38), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n602), .B(new_n603), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n599), .A2(new_n600), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n556), .A2(new_n558), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n585), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n661), .B(KEYINPUT39), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n646), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT40), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n380), .A2(new_n432), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n188), .A3(new_n651), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n674), .A2(new_n677), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n224), .ZN(G45));
  NAND3_X1  g497(.A1(new_n620), .A2(new_n380), .A3(new_n661), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT83), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n299), .A2(KEYINPUT83), .A3(new_n296), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n302), .B1(new_n690), .B2(new_n273), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n303), .B(new_n272), .C1(new_n688), .C2(new_n689), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n187), .B(new_n685), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n666), .A2(new_n695), .A3(new_n187), .A4(new_n685), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n658), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT101), .B(G146), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G48));
  INV_X1    g513(.A(new_n539), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n669), .B2(new_n590), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n189), .B1(new_n495), .B2(new_n500), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G469), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n501), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n540), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n624), .A2(new_n630), .A3(new_n701), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND3_X1  g523(.A1(new_n306), .A2(new_n609), .A3(new_n641), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n606), .A2(new_n539), .A3(new_n706), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n384), .ZN(G18));
  NAND2_X1  g527(.A1(new_n306), .A2(new_n706), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n606), .A2(new_n442), .A3(new_n651), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n207), .ZN(G21));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n679), .B(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n703), .A2(new_n609), .A3(new_n540), .A4(new_n501), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n569), .B1(new_n559), .B2(new_n565), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n595), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n592), .B1(new_n601), .B2(new_n722), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n627), .A2(new_n700), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n306), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  AOI211_X1 g540(.A(new_n188), .B(new_n705), .C1(new_n304), .C2(new_n305), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n684), .A2(KEYINPUT103), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n620), .A2(new_n380), .A3(new_n729), .A4(new_n661), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n601), .A2(new_n722), .ZN(new_n732));
  AOI21_X1  g546(.A(G902), .B1(new_n596), .B2(new_n601), .ZN(new_n733));
  OAI221_X1 g547(.A(new_n651), .B1(new_n732), .B2(new_n592), .C1(new_n625), .C2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT104), .B(G125), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G27));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n504), .B2(new_n505), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT105), .B1(new_n503), .B2(new_n493), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n741), .A2(new_n443), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n501), .A2(new_n502), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n742), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n504), .A2(new_n505), .ZN(new_n747));
  OAI211_X1 g561(.A(G469), .B(new_n746), .C1(new_n747), .C2(new_n740), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n501), .A2(new_n502), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n540), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n188), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n304), .A2(new_n751), .A3(new_n305), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n731), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n701), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n606), .A2(new_n539), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n304), .A2(new_n751), .A3(new_n305), .A4(new_n753), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  INV_X1    g578(.A(new_n662), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n754), .A2(new_n701), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n768), .A3(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND3_X1  g585(.A1(new_n304), .A2(new_n187), .A3(new_n305), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n378), .B1(new_n637), .B2(new_n361), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n620), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT110), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT43), .Z(new_n776));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n775), .B(KEYINPUT43), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  INV_X1    g594(.A(new_n651), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n645), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n772), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT44), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(G469), .B1(new_n747), .B2(KEYINPUT45), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT108), .B(G469), .C1(new_n747), .C2(KEYINPUT45), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT45), .B(new_n746), .C1(new_n747), .C2(new_n740), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n502), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n502), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n501), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n540), .A3(new_n675), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT109), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n783), .A2(new_n784), .ZN(new_n803));
  INV_X1    g617(.A(new_n772), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(KEYINPUT112), .A3(new_n786), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n789), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n540), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT47), .Z(new_n809));
  NOR4_X1   g623(.A1(new_n772), .A2(new_n606), .A3(new_n539), .A4(new_n684), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n658), .A2(new_n663), .B1(new_n727), .B2(new_n735), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n661), .A2(KEYINPUT116), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n661), .A2(KEYINPUT116), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n816), .A2(new_n817), .A3(new_n752), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n751), .A2(new_n781), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n306), .A3(new_n674), .A4(new_n719), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n815), .A2(new_n697), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n815), .A2(new_n697), .A3(KEYINPUT52), .A4(new_n820), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n825), .B1(new_n821), .B2(new_n822), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n187), .B(new_n442), .C1(new_n691), .C2(new_n692), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n652), .A2(new_n645), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n606), .A2(new_n542), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n712), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n421), .A2(new_n422), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n430), .B1(new_n429), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n423), .A2(new_n382), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n425), .A2(new_n841), .A3(new_n431), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n842), .A3(new_n372), .A4(new_n379), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n627), .A2(new_n541), .A3(new_n843), .A4(new_n602), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n666), .A3(new_n187), .A4(new_n609), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n725), .B(new_n845), .C1(new_n714), .C2(new_n715), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n623), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n306), .A2(KEYINPUT113), .A3(new_n609), .A4(new_n622), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n628), .A3(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n707), .A2(new_n836), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n842), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n639), .A2(new_n661), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n304), .A2(new_n187), .A3(new_n854), .A4(new_n305), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n627), .A2(new_n723), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n651), .A3(new_n728), .A4(new_n730), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n657), .A2(new_n855), .B1(new_n857), .B2(new_n760), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n768), .B1(new_n761), .B2(new_n765), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n759), .A2(new_n760), .A3(KEYINPUT107), .A4(new_n662), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT115), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n770), .A2(new_n864), .A3(new_n859), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n852), .A2(new_n763), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n814), .B1(new_n831), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n607), .B(new_n653), .C1(new_n710), .C2(new_n711), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n846), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n707), .A3(new_n763), .A4(new_n851), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n864), .B1(new_n770), .B2(new_n859), .ZN(new_n871));
  AOI211_X1 g685(.A(KEYINPUT115), .B(new_n858), .C1(new_n767), .C2(new_n769), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n821), .A2(new_n823), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n827), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n813), .B1(new_n867), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT53), .B1(new_n831), .B2(new_n866), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n814), .A3(new_n875), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT54), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT119), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n875), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n821), .A2(new_n822), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n824), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n826), .A3(new_n828), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n873), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n814), .B1(new_n873), .B2(new_n885), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n871), .A2(new_n872), .ZN(new_n889));
  INV_X1    g703(.A(new_n870), .ZN(new_n890));
  AND4_X1   g704(.A1(new_n814), .A2(new_n889), .A3(new_n890), .A4(new_n875), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n813), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n437), .A2(new_n779), .A3(new_n539), .A4(new_n856), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n188), .A3(new_n668), .A4(new_n706), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT50), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n779), .A2(new_n437), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n304), .A2(new_n305), .A3(new_n704), .A4(new_n753), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n734), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT120), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n704), .A2(new_n752), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n804), .B(new_n895), .C1(new_n809), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n669), .A2(new_n539), .A3(new_n673), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n905), .A2(new_n900), .A3(new_n436), .ZN(new_n906));
  INV_X1    g720(.A(new_n620), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n773), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n898), .A2(new_n902), .A3(new_n904), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT51), .ZN(new_n910));
  INV_X1    g724(.A(new_n908), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n897), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n902), .A4(new_n904), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n899), .A2(new_n759), .A3(new_n900), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT48), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n895), .A2(new_n727), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n622), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n434), .A3(new_n918), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT121), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT121), .B1(new_n916), .B2(new_n919), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n910), .A2(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n881), .A2(new_n894), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n433), .A2(new_n322), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n704), .B(KEYINPUT49), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n773), .A2(new_n620), .A3(new_n753), .ZN(new_n927));
  OR4_X1    g741(.A1(new_n667), .A2(new_n905), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(G75));
  NAND4_X1  g743(.A1(new_n878), .A2(G210), .A3(G902), .A4(new_n879), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n299), .B(new_n296), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT55), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n932), .A2(KEYINPUT122), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n322), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n932), .B2(new_n934), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT122), .B1(new_n932), .B2(new_n934), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n935), .A2(new_n938), .A3(new_n939), .ZN(G51));
  XOR2_X1   g754(.A(new_n502), .B(KEYINPUT57), .Z(new_n941));
  NOR3_X1   g755(.A1(new_n888), .A2(new_n891), .A3(new_n813), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n880), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n500), .B2(new_n495), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n888), .A2(new_n891), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(G902), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(new_n795), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n936), .B1(new_n944), .B2(new_n947), .ZN(G54));
  INV_X1    g762(.A(new_n635), .ZN(new_n949));
  NAND2_X1  g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n937), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(G60));
  NAND2_X1  g768(.A1(new_n611), .A2(new_n612), .ZN(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n615), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n955), .B(new_n957), .C1(new_n942), .C2(new_n880), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n937), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n893), .B1(new_n887), .B2(new_n892), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n955), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n888), .A2(new_n891), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n649), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n968), .B(new_n937), .C1(new_n536), .C2(new_n967), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n967), .A2(new_n536), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n937), .A3(new_n968), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G66));
  OAI21_X1  g789(.A(G953), .B1(new_n440), .B2(new_n241), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT125), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n852), .B2(G953), .ZN(new_n978));
  INV_X1    g792(.A(new_n299), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(G898), .B2(new_n322), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  AND2_X1   g795(.A1(new_n621), .A2(new_n843), .ZN(new_n982));
  NOR4_X1   g796(.A1(new_n759), .A2(new_n772), .A3(new_n676), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n809), .B2(new_n810), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n805), .A2(new_n802), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT112), .B1(new_n785), .B2(new_n786), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n815), .A2(new_n697), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n682), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT62), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n322), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n581), .A2(new_n582), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n367), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n802), .A2(new_n306), .A3(new_n701), .A4(new_n719), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n994), .A2(new_n811), .A3(new_n763), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n988), .B1(new_n769), .B2(new_n767), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n806), .A2(new_n995), .A3(new_n322), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(G900), .B2(G953), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n991), .A2(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT126), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1001), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1000), .B1(new_n999), .B2(new_n1002), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  OR2_X1    g823(.A1(new_n987), .A2(new_n990), .ZN(new_n1010));
  INV_X1    g824(.A(new_n852), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n584), .A3(new_n569), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n806), .A2(new_n995), .A3(new_n996), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1009), .B1(new_n1014), .B2(new_n1011), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n555), .A3(new_n583), .A4(new_n585), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n599), .A2(new_n600), .A3(new_n586), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1009), .B(new_n1017), .C1(new_n882), .C2(new_n886), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n937), .A2(new_n1013), .A3(new_n1016), .A4(new_n1018), .ZN(G57));
endmodule


