//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n204), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT66), .B(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n221), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT67), .Z(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G116), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n209), .A2(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n251), .A2(new_n255), .A3(new_n217), .A4(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n254), .B1(new_n257), .B2(new_n253), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n217), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT86), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT86), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n259), .A2(new_n263), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G283), .ZN(new_n265));
  INV_X1    g0065(.A(G97), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n265), .B(new_n210), .C1(G33), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n262), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  XOR2_X1   g0068(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n269));
  AOI21_X1  g0069(.A(new_n258), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n262), .A2(new_n271), .A3(new_n264), .A4(new_n267), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G264), .A3(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G257), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G303), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n275), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT5), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT81), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(G1), .A2(G13), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(G270), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n291), .B2(new_n292), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(new_n287), .A3(new_n285), .A4(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT84), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n294), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n282), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT85), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT85), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n282), .B(new_n303), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(G200), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n302), .A2(new_n304), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n274), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n270), .B2(new_n272), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT21), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n302), .A2(KEYINPUT21), .A3(new_n304), .A4(new_n310), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n282), .B(G179), .C1(new_n299), .C2(new_n300), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n273), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n308), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n210), .A2(G33), .ZN(new_n321));
  INV_X1    g0121(.A(G150), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G20), .A2(G33), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n320), .A2(new_n321), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n259), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n252), .A2(new_n259), .ZN(new_n328));
  INV_X1    g0128(.A(G50), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n209), .B2(G20), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(new_n330), .B1(new_n329), .B2(new_n252), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT9), .ZN(new_n333));
  AOI21_X1  g0133(.A(G1), .B1(new_n286), .B2(new_n288), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n293), .A2(G274), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n293), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G222), .A2(G1698), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n277), .A2(G223), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n275), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n281), .C1(G77), .C2(new_n275), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(G190), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G200), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n333), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT10), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n309), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n340), .A2(new_n353), .A3(new_n344), .A4(new_n345), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n332), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT70), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n259), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n251), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n209), .A2(G20), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G77), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n359), .A2(new_n361), .B1(G77), .B2(new_n251), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G20), .A2(G77), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n363), .B1(new_n364), .B2(new_n321), .C1(new_n324), .C2(new_n320), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n259), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G244), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n335), .B1(new_n337), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n275), .A2(G232), .A3(new_n277), .ZN(new_n370));
  INV_X1    g0170(.A(G107), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n275), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n372), .B2(new_n281), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n366), .B1(new_n374), .B2(new_n309), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n353), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n366), .B(KEYINPUT71), .C1(new_n373), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(G190), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n366), .B1(new_n373), .B2(new_n379), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n351), .A2(new_n357), .A3(new_n378), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G33), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G33), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(G223), .A4(new_n277), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT76), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n275), .A2(new_n394), .A3(G223), .A4(new_n277), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n389), .A2(new_n391), .A3(G226), .A4(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n293), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G232), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n335), .B1(new_n337), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n403), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n399), .B1(new_n395), .B2(new_n393), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(G190), .C1(new_n406), .C2(new_n293), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n324), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G58), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n204), .B1(new_n222), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n411), .B1(new_n413), .B2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n389), .A2(new_n391), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n390), .A2(G33), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT74), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n275), .B2(G20), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n222), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT75), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n414), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n210), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n419), .B1(new_n417), .B2(KEYINPUT74), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n422), .A2(new_n428), .B1(new_n429), .B2(new_n416), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n430), .A2(KEYINPUT75), .A3(new_n222), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n409), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G68), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT66), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT66), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G68), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n203), .B1(new_n437), .B2(G58), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n438), .A2(new_n210), .B1(new_n410), .B2(new_n324), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n389), .A2(new_n391), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n420), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n433), .B1(new_n423), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n358), .B1(new_n443), .B2(KEYINPUT16), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n432), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n320), .B1(new_n209), .B2(G20), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n328), .B1(new_n252), .B2(new_n320), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n408), .A2(new_n445), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n448), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n432), .B2(new_n444), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(new_n446), .A3(KEYINPUT17), .A4(new_n408), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(new_n448), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  OAI21_X1  g0257(.A(G169), .B1(new_n401), .B2(new_n403), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n405), .B(G179), .C1(new_n406), .C2(new_n293), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT18), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  INV_X1    g0262(.A(new_n460), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n453), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT7), .B1(new_n440), .B2(new_n210), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n275), .A2(new_n419), .ZN(new_n467));
  OAI21_X1  g0267(.A(G68), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n259), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT75), .B1(new_n430), .B2(new_n222), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n424), .A2(new_n425), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n414), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n473), .B2(new_n409), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT18), .B(new_n460), .C1(new_n474), .C2(new_n452), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT77), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n455), .B1(new_n465), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n437), .A2(new_n210), .ZN(new_n478));
  INV_X1    g0278(.A(G77), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n324), .A2(new_n329), .B1(new_n321), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n259), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n482), .A2(KEYINPUT11), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(KEYINPUT11), .ZN(new_n484));
  INV_X1    g0284(.A(G13), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n478), .A2(KEYINPUT12), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n328), .A2(G68), .A3(new_n360), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n251), .A2(G68), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(KEYINPUT12), .C2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n483), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT14), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n335), .B1(new_n337), .B2(new_n223), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n338), .A2(new_n277), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n402), .A2(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n389), .A2(new_n494), .A3(new_n391), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n293), .B1(new_n498), .B2(KEYINPUT72), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT72), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  AOI211_X1 g0301(.A(KEYINPUT13), .B(new_n493), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT13), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(KEYINPUT72), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n281), .A3(new_n501), .ZN(new_n505));
  INV_X1    g0305(.A(new_n493), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n492), .B(G169), .C1(new_n502), .C2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n496), .A2(new_n500), .A3(new_n497), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n500), .B1(new_n496), .B2(new_n497), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n509), .A2(new_n510), .A3(new_n293), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT13), .B1(new_n511), .B2(new_n493), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n503), .A3(new_n506), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(G179), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n492), .B1(new_n516), .B2(G169), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT73), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(G169), .B1(new_n502), .B2(new_n507), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT73), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n514), .A4(new_n508), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n491), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(G200), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n512), .A2(G190), .A3(new_n513), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n491), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n387), .A2(new_n477), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n290), .A2(new_n293), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n389), .A2(new_n391), .A3(G257), .A4(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n389), .A2(new_n391), .A3(G250), .A4(new_n277), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G294), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n531), .A2(G264), .B1(new_n535), .B2(new_n281), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(KEYINPUT88), .A3(new_n307), .A4(new_n297), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT88), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n281), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n290), .A2(G264), .A3(new_n293), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n297), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n379), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(G190), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n257), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n371), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT25), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n251), .B2(G107), .ZN(new_n548));
  AOI22_X1  g0348(.A1(G107), .A2(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n389), .A2(new_n391), .A3(new_n210), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n275), .A2(new_n553), .A3(new_n210), .A4(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(G20), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n210), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n371), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT24), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n555), .A2(new_n564), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n550), .B1(new_n566), .B2(new_n259), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n544), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n555), .A2(new_n564), .A3(new_n561), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n564), .B1(new_n555), .B2(new_n561), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n259), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n549), .ZN(new_n572));
  INV_X1    g0372(.A(new_n541), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n353), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n541), .A2(new_n309), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT89), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n568), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n371), .B1(new_n421), .B2(new_n423), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n324), .A2(new_n479), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n371), .A2(KEYINPUT6), .A3(G97), .ZN(new_n585));
  XNOR2_X1  g0385(.A(G97), .B(G107), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT6), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n584), .B1(new_n588), .B2(new_n210), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n259), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n251), .A2(G97), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n545), .B2(G97), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G257), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n297), .B1(new_n530), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n389), .A2(new_n391), .A3(G244), .A4(new_n277), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT79), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT79), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n389), .A2(new_n391), .A3(G250), .A4(G1698), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n603), .A2(new_n265), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n595), .B1(new_n605), .B2(new_n281), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n593), .B1(G190), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT80), .ZN(new_n608));
  INV_X1    g0408(.A(new_n601), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n265), .B(new_n603), .C1(new_n596), .C2(new_n597), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n600), .B1(new_n596), .B2(new_n597), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n608), .B1(new_n612), .B2(new_n293), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n605), .A2(KEYINPUT80), .A3(new_n281), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n595), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n607), .B1(new_n615), .B2(new_n379), .ZN(new_n616));
  INV_X1    g0416(.A(new_n595), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n605), .A2(KEYINPUT80), .A3(new_n281), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT80), .B1(new_n605), .B2(new_n281), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n353), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n592), .ZN(new_n621));
  AND2_X1   g0421(.A1(G97), .A2(G107), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n587), .B1(new_n622), .B2(new_n206), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n371), .A2(KEYINPUT6), .A3(G97), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n583), .B1(new_n625), .B2(G20), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n430), .B2(new_n371), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n621), .B1(new_n627), .B2(new_n259), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n617), .B1(new_n612), .B2(new_n293), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n309), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(G250), .B1(new_n288), .B2(G1), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n281), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n293), .A2(G274), .A3(new_n289), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT82), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT82), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n296), .A2(new_n636), .A3(new_n289), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n389), .A2(new_n391), .A3(G244), .A4(G1698), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n556), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT83), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n275), .A2(new_n641), .A3(G238), .A4(new_n277), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n389), .A2(new_n391), .A3(G238), .A4(new_n277), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT83), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n638), .B(new_n353), .C1(new_n645), .C2(new_n293), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT19), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n210), .B1(new_n497), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(G87), .B2(new_n207), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n389), .A2(new_n391), .A3(new_n210), .A4(G68), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n647), .B1(new_n321), .B2(new_n266), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n259), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n364), .A2(new_n252), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(new_n257), .C2(new_n364), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n638), .B1(new_n645), .B2(new_n293), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n309), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n545), .A2(G87), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n653), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n657), .B2(G200), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n638), .B(G190), .C1(new_n645), .C2(new_n293), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n656), .A2(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n616), .A2(new_n631), .A3(new_n663), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n319), .A2(new_n529), .A3(new_n581), .A4(new_n664), .ZN(G372));
  AND2_X1   g0465(.A1(new_n451), .A2(new_n454), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n527), .A2(new_n377), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n523), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n464), .A2(new_n475), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n351), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n357), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n387), .A2(new_n528), .A3(new_n477), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n658), .A2(new_n646), .A3(new_n655), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n593), .B1(new_n606), .B2(G169), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n615), .B2(new_n353), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT26), .B1(new_n676), .B2(new_n663), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n657), .A2(G200), .ZN(new_n678));
  INV_X1    g0478(.A(new_n660), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n662), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n631), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n674), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  AND4_X1   g0484(.A1(new_n313), .A2(new_n317), .A3(new_n314), .A4(new_n576), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n616), .A2(new_n631), .A3(new_n568), .A4(new_n663), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n672), .B1(new_n673), .B2(new_n688), .ZN(G369));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n486), .A2(new_n210), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT90), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G213), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n691), .B2(KEYINPUT27), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n273), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n318), .A2(new_n313), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n319), .A2(KEYINPUT93), .ZN(new_n705));
  INV_X1    g0505(.A(new_n701), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n319), .A2(KEYINPUT93), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n690), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n699), .A2(new_n572), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n581), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT94), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n581), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  INV_X1    g0514(.A(new_n576), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n712), .A2(new_n714), .B1(new_n715), .B2(new_n699), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n698), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n699), .B1(new_n318), .B2(new_n313), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n712), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n213), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(G87), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n206), .A2(new_n725), .A3(new_n253), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT95), .Z(new_n727));
  NOR3_X1   g0527(.A1(new_n724), .A2(new_n727), .A3(new_n209), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n220), .B2(new_n724), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  OAI21_X1  g0530(.A(new_n698), .B1(new_n684), .B2(new_n687), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G200), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n734), .A2(new_n607), .B1(new_n620), .B2(new_n630), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n313), .A2(new_n317), .A3(new_n576), .A4(new_n314), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n568), .A4(new_n663), .ZN(new_n737));
  INV_X1    g0537(.A(new_n674), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n620), .A2(new_n630), .A3(new_n674), .A4(new_n680), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n682), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n663), .A2(KEYINPUT26), .A3(new_n620), .A4(new_n630), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n699), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n732), .A2(new_n745), .ZN(new_n746));
  AND4_X1   g0546(.A1(new_n319), .A2(new_n581), .A3(new_n664), .A4(new_n698), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n644), .A2(new_n642), .ZN(new_n748));
  INV_X1    g0548(.A(new_n640), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n293), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n635), .A2(new_n637), .ZN(new_n751));
  INV_X1    g0551(.A(new_n633), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n754), .A2(new_n573), .A3(G179), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n306), .A2(new_n733), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n606), .A2(new_n754), .A3(new_n536), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(new_n315), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n539), .A2(new_n540), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n657), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n316), .A2(new_n761), .A3(KEYINPUT30), .A4(new_n606), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n699), .B1(new_n756), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n306), .A2(new_n733), .A3(new_n755), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n759), .A3(new_n762), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(G330), .B1(new_n747), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n746), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n730), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(new_n485), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n209), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n724), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n709), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n704), .A2(new_n708), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(G330), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  INV_X1    g0582(.A(new_n778), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n213), .A2(G355), .A3(new_n275), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n723), .A2(new_n275), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n219), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n246), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n784), .B(new_n787), .C1(new_n253), .C2(new_n723), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n217), .B1(G20), .B2(new_n309), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n783), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n210), .A2(new_n307), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n353), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n210), .A2(G190), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G58), .A2(new_n800), .B1(new_n803), .B2(G77), .ZN(new_n804));
  NAND3_X1  g0604(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n307), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n804), .B1(new_n329), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT97), .Z(new_n809));
  NOR2_X1   g0609(.A1(G179), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n801), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G159), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n805), .A2(G190), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n210), .B1(new_n810), .B2(G190), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n433), .B1(new_n817), .B2(new_n266), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n379), .A2(G179), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n801), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n371), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n797), .A2(new_n819), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n275), .B1(new_n822), .B2(new_n725), .ZN(new_n823));
  NOR4_X1   g0623(.A1(new_n814), .A2(new_n818), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G322), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n799), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n827), .A2(new_n820), .B1(new_n802), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n829), .C1(G329), .C2(new_n812), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n440), .B1(new_n822), .B2(new_n279), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT33), .B(G317), .Z(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n816), .A2(new_n832), .B1(new_n833), .B2(new_n817), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n834), .C1(G326), .C2(new_n806), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n809), .A2(new_n824), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n792), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n795), .B1(new_n796), .B2(new_n836), .C1(new_n780), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n782), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n377), .A2(new_n699), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n698), .A2(new_n366), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n382), .B2(new_n385), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n378), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n731), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n698), .B(new_n848), .C1(new_n684), .C2(new_n687), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n778), .B1(new_n850), .B2(new_n771), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n771), .B2(new_n850), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n796), .A2(new_n791), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n778), .B1(G77), .B2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT98), .Z(new_n855));
  OAI221_X1 g0655(.A(new_n440), .B1(new_n817), .B2(new_n266), .C1(new_n833), .C2(new_n799), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n816), .A2(new_n827), .B1(new_n807), .B2(new_n279), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n822), .A2(new_n371), .B1(new_n820), .B2(new_n725), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n802), .A2(new_n253), .B1(new_n811), .B2(new_n828), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n800), .B1(new_n803), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n861), .B1(new_n807), .B2(new_n862), .C1(new_n322), .C2(new_n816), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT34), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n817), .A2(new_n412), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n275), .B1(new_n822), .B2(new_n329), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n820), .A2(new_n433), .B1(new_n811), .B2(new_n868), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n863), .A2(new_n864), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n855), .B1(new_n796), .B2(new_n872), .C1(new_n848), .C2(new_n791), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n852), .A2(new_n873), .ZN(G384));
  NOR2_X1   g0674(.A1(new_n775), .A2(new_n209), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n443), .A2(KEYINPUT16), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n448), .B1(new_n876), .B2(new_n470), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n697), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n476), .A2(new_n461), .A3(new_n464), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(new_n455), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n453), .A2(new_n408), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n877), .B1(new_n460), .B2(new_n697), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n460), .B1(new_n474), .B2(new_n452), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n697), .B1(new_n474), .B2(new_n452), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n882), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n887), .B1(new_n666), .B2(new_n669), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n886), .A2(new_n887), .A3(new_n882), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(new_n889), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n892), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n518), .A2(new_n522), .ZN(new_n900));
  INV_X1    g0700(.A(new_n491), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n491), .A2(new_n698), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n526), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n523), .B2(new_n527), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n846), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n768), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT31), .B1(new_n768), .B2(new_n699), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n319), .A2(new_n581), .A3(new_n664), .A4(new_n698), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n899), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n881), .B2(new_n890), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n476), .A2(new_n461), .A3(new_n464), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n878), .B1(new_n666), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n890), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n917), .A2(new_n918), .A3(new_n892), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n912), .B(new_n907), .C1(new_n915), .C2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(KEYINPUT102), .A3(new_n921), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n914), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT103), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n529), .A2(new_n912), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n690), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n927), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n892), .B1(new_n917), .B2(new_n918), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n891), .A2(new_n932), .A3(KEYINPUT39), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT39), .B1(new_n891), .B2(new_n897), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n902), .A2(new_n699), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n669), .A2(new_n697), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n891), .A2(new_n932), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n842), .B(KEYINPUT100), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n849), .A2(new_n941), .B1(new_n905), .B2(new_n906), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n529), .B1(new_n732), .B2(new_n745), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n945), .A2(new_n672), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n944), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n875), .B1(new_n931), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n931), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n220), .B(G77), .C1(new_n412), .C2(new_n222), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n433), .B2(new_n202), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(G1), .A3(new_n485), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(G116), .A4(new_n218), .ZN(new_n956));
  XNOR2_X1  g0756(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n950), .A2(new_n953), .A3(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT104), .Z(G367));
  OAI21_X1  g0760(.A(new_n794), .B1(new_n213), .B2(new_n364), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n785), .B2(new_n242), .ZN(new_n962));
  INV_X1    g0762(.A(new_n822), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(G116), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n802), .A2(new_n827), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n820), .A2(new_n266), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(G317), .C2(new_n812), .ZN(new_n968));
  INV_X1    g0768(.A(new_n817), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n969), .A2(G107), .B1(G311), .B2(new_n806), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n440), .B1(new_n799), .B2(new_n279), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G294), .B2(new_n815), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n965), .A2(new_n968), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n275), .B1(new_n802), .B2(new_n201), .C1(new_n816), .C2(new_n410), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G143), .B2(new_n806), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n822), .A2(new_n412), .B1(new_n820), .B2(new_n479), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G137), .B2(new_n812), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n969), .A2(G68), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n322), .B2(new_n799), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT107), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n973), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT47), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n783), .B(new_n962), .C1(new_n983), .C2(new_n793), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n698), .A2(new_n679), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n738), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n681), .B2(new_n985), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n984), .B1(new_n837), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n724), .B(KEYINPUT41), .Z(new_n989));
  OAI21_X1  g0789(.A(new_n735), .B1(new_n628), .B2(new_n698), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n676), .A2(new_n699), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n721), .A2(new_n719), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n992), .B1(new_n721), .B2(new_n719), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT44), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n997), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n718), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(KEYINPUT106), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n997), .B(new_n718), .C1(new_n999), .C2(new_n1001), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT106), .B1(new_n709), .B2(new_n717), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n720), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n716), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n721), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n709), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n709), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n721), .A3(new_n1008), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n772), .B(new_n1006), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1004), .A2(new_n1005), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n989), .B1(new_n1015), .B2(new_n773), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n777), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n992), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n718), .A2(KEYINPUT105), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT105), .B1(new_n718), .B2(new_n1018), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n715), .A2(new_n616), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n699), .B1(new_n1024), .B2(new_n631), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1010), .A2(new_n992), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT42), .B2(new_n1026), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1020), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1023), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1030), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n988), .B1(new_n1017), .B2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n773), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1011), .A2(new_n1013), .A3(new_n772), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n724), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n716), .A2(new_n792), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n822), .A2(new_n833), .B1(new_n817), .B2(new_n827), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G317), .A2(new_n800), .B1(new_n803), .B2(G303), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n807), .B2(new_n825), .C1(new_n828), .C2(new_n816), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n820), .A2(new_n253), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n275), .B(new_n1050), .C1(G326), .C2(new_n812), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n440), .B(new_n967), .C1(G159), .C2(new_n806), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G68), .A2(new_n803), .B1(new_n812), .B2(G150), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G50), .A2(new_n800), .B1(new_n963), .B2(G77), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n364), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n320), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1056), .A2(new_n969), .B1(new_n1057), .B2(new_n815), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n796), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n785), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n239), .B2(G45), .ZN(new_n1062));
  AOI211_X1 g0862(.A(G45), .B(new_n727), .C1(G68), .C2(G77), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT108), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n320), .A2(G50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1062), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n727), .A2(new_n213), .A3(new_n275), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G107), .C2(new_n213), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n783), .B(new_n1060), .C1(new_n794), .C2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1036), .A2(new_n777), .B1(new_n1040), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1039), .A2(new_n1073), .ZN(G393));
  OAI221_X1 g0874(.A(new_n794), .B1(new_n266), .B2(new_n213), .C1(new_n1061), .C2(new_n249), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(new_n778), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n807), .A2(new_n322), .B1(new_n799), .B2(new_n410), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n820), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n440), .B1(new_n1079), .B2(G87), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n437), .A2(new_n963), .B1(new_n812), .B2(G143), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n817), .A2(new_n479), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1057), .B2(new_n803), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n201), .B2(new_n816), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT109), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n800), .A2(G311), .B1(G317), .B2(new_n806), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n822), .A2(new_n827), .B1(new_n811), .B2(new_n825), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1088), .A2(new_n275), .A3(new_n821), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n802), .A2(new_n833), .B1(new_n817), .B2(new_n253), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G303), .B2(new_n815), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT110), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1082), .A2(new_n1086), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1076), .B1(new_n796), .B2(new_n1094), .C1(new_n992), .C2(new_n837), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1005), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1097), .B2(new_n776), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1015), .A2(new_n724), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1037), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(new_n724), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n690), .B1(new_n910), .B2(new_n911), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n907), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT39), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n669), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n456), .B(new_n697), .C1(new_n1108), .C2(new_n455), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n895), .A2(new_n889), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT38), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1107), .B1(new_n919), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n891), .A2(new_n932), .A3(KEYINPUT39), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n905), .A2(new_n906), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n699), .B(new_n846), .C1(new_n737), .C2(new_n742), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n940), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n936), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1112), .A2(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n919), .A2(new_n1111), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1119), .A2(new_n942), .A3(new_n936), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1106), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n940), .B1(new_n743), .B2(new_n848), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n904), .B1(new_n902), .B2(new_n526), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n523), .A2(new_n527), .A3(new_n903), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1117), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n933), .B2(new_n934), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1116), .A2(new_n898), .A3(new_n1117), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1105), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1114), .B1(new_n1104), .B2(new_n848), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1122), .B1(new_n1106), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(G330), .B(new_n848), .C1(new_n747), .C2(new_n770), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1125), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1122), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1105), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT111), .B1(new_n771), .B2(new_n673), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT111), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1104), .A2(new_n529), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1132), .A2(new_n946), .A3(new_n1136), .A4(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1130), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1103), .B1(new_n1142), .B2(KEYINPUT113), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT112), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n771), .A2(KEYINPUT111), .A3(new_n673), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1138), .B1(new_n1104), .B2(new_n529), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n672), .B(new_n945), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1134), .A2(new_n1135), .A3(new_n1105), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1135), .B1(new_n1134), .B2(new_n1105), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT112), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n1121), .A4(new_n1129), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1144), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1143), .B(new_n1153), .C1(KEYINPUT113), .C2(new_n1142), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n778), .B1(new_n1057), .B2(new_n853), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n935), .A2(new_n791), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n275), .B1(new_n820), .B2(new_n201), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT115), .Z(new_n1158));
  NOR2_X1   g0958(.A1(new_n822), .A2(new_n322), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT53), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n802), .A2(new_n1161), .B1(new_n811), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G132), .B2(new_n800), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1158), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n969), .A2(G159), .B1(G128), .B2(new_n806), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n862), .B2(new_n816), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1083), .B1(new_n815), .B2(G107), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n827), .B2(new_n807), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n820), .A2(new_n433), .B1(new_n811), .B2(new_n833), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT116), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT116), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n275), .B1(new_n963), .B2(G87), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G116), .A2(new_n800), .B1(new_n803), .B2(G97), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1165), .A2(new_n1167), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1155), .B(new_n1156), .C1(new_n793), .C2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1130), .A2(new_n776), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1178), .A2(KEYINPUT114), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(KEYINPUT114), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1154), .A2(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n671), .A2(new_n355), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n697), .A2(new_n332), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1185), .B(new_n1186), .Z(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n926), .B2(G330), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n899), .A2(new_n913), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n920), .A2(KEYINPUT102), .A3(new_n921), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT102), .B1(new_n920), .B2(new_n921), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n1190), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n1187), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n944), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n926), .A2(G330), .A3(new_n1188), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1187), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n944), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1147), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1195), .A2(new_n1199), .B1(new_n1153), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n724), .B1(new_n1201), .B2(KEYINPUT57), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT119), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1195), .A2(new_n1203), .A3(new_n1199), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1153), .B2(new_n1200), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1196), .A2(new_n1197), .A3(KEYINPUT119), .A4(new_n1198), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1187), .A2(new_n790), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n778), .B1(new_n202), .B2(new_n853), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n275), .A2(G41), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G50), .B(new_n1213), .C1(new_n388), .C2(new_n286), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n979), .B(new_n1213), .C1(new_n479), .C2(new_n822), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n364), .A2(new_n802), .B1(new_n820), .B2(new_n412), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n816), .A2(new_n266), .B1(new_n807), .B2(new_n253), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n799), .A2(new_n371), .B1(new_n811), .B2(new_n827), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1220));
  AOI21_X1  g1020(.A(new_n1214), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n969), .A2(G150), .B1(G125), .B2(new_n806), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT118), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n816), .A2(new_n868), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n800), .A2(G128), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n822), .A2(new_n1161), .B1(new_n802), .B2(new_n862), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT59), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n388), .B(new_n286), .C1(new_n820), .C2(new_n410), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G124), .B2(new_n812), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .C1(new_n1229), .C2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1212), .B1(new_n1233), .B2(new_n793), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1210), .A2(new_n777), .B1(new_n1211), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1209), .A2(new_n1235), .ZN(G375));
  NOR3_X1   g1036(.A1(new_n1148), .A2(new_n1149), .A3(new_n776), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1125), .A2(new_n790), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n778), .B1(G68), .B2(new_n853), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n822), .A2(new_n266), .B1(new_n811), .B2(new_n279), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT120), .Z(new_n1241));
  AOI22_X1  g1041(.A1(G283), .A2(new_n800), .B1(new_n803), .B2(G107), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n275), .B1(new_n1079), .B2(G77), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n806), .A2(G294), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n969), .A2(new_n1056), .B1(G116), .B2(new_n815), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n440), .B1(new_n1079), .B2(G58), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n329), .B2(new_n817), .C1(new_n816), .C2(new_n1161), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G159), .A2(new_n963), .B1(new_n803), .B2(G150), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G137), .A2(new_n800), .B1(new_n812), .B2(G128), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n806), .A2(KEYINPUT121), .A3(G132), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n807), .B2(new_n868), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1241), .A2(new_n1246), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1239), .B1(new_n1255), .B2(new_n793), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1237), .B1(new_n1238), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n989), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1141), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G381));
  NOR2_X1   g1061(.A1(G396), .A2(G393), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G378), .A2(new_n1263), .A3(G384), .A4(G381), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1032), .B(new_n1033), .C1(new_n1016), .C2(new_n777), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1265), .A2(new_n988), .A3(new_n1101), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1209), .A3(new_n1235), .A4(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n695), .A2(G343), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT122), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(G375), .C2(new_n1271), .ZN(G409));
  XNOR2_X1  g1072(.A(G393), .B(new_n840), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1101), .B1(new_n1265), .B2(new_n988), .ZN(new_n1274));
  OAI211_X1 g1074(.A(KEYINPUT123), .B(new_n1273), .C1(new_n1266), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(G390), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1273), .A2(KEYINPUT123), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1265), .A2(new_n1101), .A3(new_n988), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(KEYINPUT123), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1275), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1235), .C1(new_n1202), .C2(new_n1208), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1204), .A2(new_n777), .A3(new_n1207), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1211), .A2(new_n1234), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1153), .A2(new_n1200), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1210), .A2(new_n1259), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1268), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1269), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1292), .A2(new_n1258), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n724), .B1(new_n1292), .B2(new_n1258), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1257), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n852), .A3(new_n873), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G384), .B(new_n1257), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G2897), .ZN(new_n1299));
  OR3_X1    g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1269), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1270), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1302), .A2(new_n1299), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1282), .B1(new_n1291), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1290), .A2(new_n1269), .A3(new_n1301), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1270), .B1(new_n1283), .B2(new_n1289), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1298), .A2(new_n1307), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1310), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1305), .B(new_n1308), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1290), .A2(new_n1302), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1304), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n1270), .B(new_n1320), .C1(new_n1283), .C2(new_n1289), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1319), .A2(new_n1321), .B1(new_n1306), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1315), .B2(new_n1320), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1318), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1275), .A2(new_n1280), .A3(KEYINPUT127), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT127), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1314), .B1(new_n1325), .B2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1268), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1283), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1301), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1283), .A3(new_n1298), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1328), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1326), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1327), .ZN(new_n1337));
  AOI22_X1  g1137(.A1(new_n1333), .A2(new_n1334), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1335), .A2(new_n1338), .ZN(G402));
endmodule


