//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n628, new_n629, new_n631, new_n632, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n451), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT70), .B(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(new_n463), .A3(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT71), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(KEYINPUT71), .A3(new_n468), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(G160));
  OAI221_X1 g047(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n473));
  INV_X1    g048(.A(G124), .ZN(new_n474));
  INV_X1    g049(.A(new_n463), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n461), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n461), .A2(new_n466), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT72), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n461), .A2(new_n480), .A3(new_n466), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n477), .B1(G136), .B2(new_n482), .ZN(G162));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(KEYINPUT73), .B2(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n461), .A2(new_n463), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n461), .A2(new_n463), .A3(new_n490), .A4(new_n485), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n466), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n461), .A2(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT74), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT75), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n506), .A3(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n500), .A2(new_n501), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n504), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n507), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n509), .B1(new_n506), .B2(G543), .ZN(new_n522));
  NOR3_X1   g097(.A1(new_n499), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n519), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI211_X1 g101(.A(G51), .B(G543), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n524), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n508), .A2(new_n510), .ZN(new_n534));
  AND4_X1   g109(.A1(G89), .A2(new_n534), .A3(new_n519), .A4(new_n512), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT76), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n511), .A2(G89), .A3(new_n512), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n532), .A2(new_n527), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n524), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(G168));
  XOR2_X1   g116(.A(KEYINPUT78), .B(G52), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n502), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n513), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n511), .A2(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n516), .B1(new_n548), .B2(KEYINPUT77), .ZN(new_n549));
  INV_X1    g124(.A(G77), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n499), .ZN(new_n551));
  AOI211_X1 g126(.A(KEYINPUT77), .B(new_n551), .C1(new_n511), .C2(G64), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n545), .B1(new_n549), .B2(new_n553), .ZN(G171));
  AND2_X1   g129(.A1(G68), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n511), .B2(G56), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n516), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n511), .A2(G81), .A3(new_n512), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n502), .A2(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND3_X1  g141(.A1(new_n511), .A2(G91), .A3(new_n512), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n525), .C2(new_n526), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OAI221_X1 g146(.A(new_n567), .B1(new_n569), .B2(new_n570), .C1(new_n571), .C2(new_n516), .ZN(G299));
  INV_X1    g147(.A(new_n513), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G90), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n551), .B1(new_n511), .B2(G64), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n574), .B(new_n543), .C1(new_n577), .C2(new_n552), .ZN(G301));
  AND3_X1   g153(.A1(new_n536), .A2(KEYINPUT79), .A3(new_n540), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT79), .B1(new_n536), .B2(new_n540), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G286));
  OAI221_X1 g157(.A(new_n504), .B1(new_n505), .B2(new_n513), .C1(new_n516), .C2(new_n515), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  INV_X1    g160(.A(new_n502), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n584), .B1(new_n585), .B2(new_n586), .C1(new_n587), .C2(new_n513), .ZN(G288));
  NAND2_X1  g163(.A1(new_n511), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n516), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n573), .A2(G86), .B1(G48), .B2(new_n502), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n502), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n513), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(new_n502), .A2(G54), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n534), .A2(G66), .A3(new_n519), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n604), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n534), .A2(G92), .A3(new_n519), .A4(new_n512), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n511), .A2(KEYINPUT10), .A3(G92), .A4(new_n512), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G171), .B2(new_n615), .ZN(G284));
  OAI21_X1  g192(.A(new_n616), .B1(G171), .B2(new_n615), .ZN(G321));
  OAI21_X1  g193(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n511), .A2(G65), .ZN(new_n620));
  NAND2_X1  g195(.A1(G78), .A2(G543), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n516), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT81), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n581), .B2(G868), .ZN(G297));
  AOI21_X1  g201(.A(new_n625), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(new_n614), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g208(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n634));
  XNOR2_X1  g209(.A(G323), .B(new_n634), .ZN(G282));
  INV_X1    g210(.A(new_n476), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G123), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n475), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  INV_X1    g217(.A(new_n482), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n637), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n461), .A2(new_n467), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT13), .ZN(new_n651));
  AOI22_X1  g226(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(G2096), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n652), .B(new_n653), .C1(new_n648), .C2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(G156));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n648), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n647), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  XOR2_X1   g269(.A(G1981), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n694), .B(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT89), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT32), .B(G1981), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT88), .B(G16), .Z(new_n709));
  MUX2_X1   g284(.A(G303), .B(G22), .S(new_n709), .Z(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT33), .B(G1976), .Z(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NAND4_X1  g293(.A1(new_n706), .A2(new_n708), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n721));
  NOR2_X1   g296(.A1(G25), .A2(G29), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT86), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n482), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n636), .A2(G119), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT87), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n722), .B1(new_n728), .B2(G29), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n601), .A2(new_n709), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G24), .B2(new_n709), .ZN(new_n734));
  INV_X1    g309(.A(G1986), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT90), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n729), .A2(new_n731), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n720), .A2(new_n721), .A3(new_n732), .A4(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n482), .A2(G139), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  AOI22_X1  g322(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n747), .C1(new_n463), .C2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  MUX2_X1   g325(.A(G33), .B(new_n750), .S(G29), .Z(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G2072), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n709), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n623), .B2(new_n713), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  INV_X1    g332(.A(G34), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(KEYINPUT24), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G160), .B2(new_n757), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n756), .B1(G2084), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT26), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n766), .A2(new_n767), .B1(G105), .B2(new_n467), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n476), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n482), .B2(G141), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n757), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n757), .B2(G32), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT31), .B(G11), .Z(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n757), .B1(new_n779), .B2(G28), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n781), .A2(KEYINPUT95), .B1(new_n779), .B2(G28), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n777), .B(new_n784), .C1(new_n757), .C2(new_n645), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n757), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n757), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G2084), .B2(new_n762), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n773), .A2(new_n776), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n785), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G171), .A2(new_n713), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G5), .B2(new_n713), .ZN(new_n794));
  INV_X1    g369(.A(G1961), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n752), .A2(new_n763), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n757), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT92), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT28), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n482), .A2(G140), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT91), .Z(new_n802));
  OR2_X1    g377(.A1(new_n463), .A2(G116), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n636), .A2(G128), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n800), .B1(new_n807), .B2(new_n757), .ZN(new_n808));
  INV_X1    g383(.A(G2067), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G21), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G168), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1966), .Z(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n813), .C1(new_n795), .C2(new_n794), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n757), .A2(G35), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G162), .B2(new_n757), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT29), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G2090), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT96), .Z(new_n819));
  NOR2_X1   g394(.A1(G4), .A2(G16), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n628), .B2(G16), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G1348), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n817), .B2(G2090), .ZN(new_n823));
  INV_X1    g398(.A(new_n561), .ZN(new_n824));
  MUX2_X1   g399(.A(new_n824), .B(G19), .S(new_n709), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1341), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(G1348), .ZN(new_n827));
  OR3_X1    g402(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n797), .A2(new_n814), .A3(new_n819), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n743), .A2(new_n744), .A3(new_n829), .ZN(G311));
  NAND3_X1  g405(.A1(new_n743), .A2(new_n744), .A3(new_n829), .ZN(G150));
  NAND2_X1  g406(.A1(new_n628), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n556), .A2(new_n516), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n511), .A2(G67), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G651), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n558), .A2(new_n559), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n511), .A2(G93), .A3(new_n512), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n502), .A2(G55), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n834), .A2(new_n838), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n516), .B1(new_n835), .B2(new_n836), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n841), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n557), .A2(new_n560), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n833), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT97), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT98), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n844), .A2(new_n845), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(G145));
  XOR2_X1   g435(.A(new_n727), .B(KEYINPUT87), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n650), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n482), .A2(G142), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n463), .A2(new_n864), .A3(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n463), .B2(G118), .ZN(new_n866));
  OR2_X1    g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n865), .A2(G2104), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n636), .A2(G130), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n728), .B(new_n650), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n771), .B(new_n497), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n807), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n749), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n875), .B(new_n878), .C1(new_n750), .C2(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n750), .B2(new_n877), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n872), .A3(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n645), .B(KEYINPUT99), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G160), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G162), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n881), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g466(.A1(new_n857), .A2(new_n615), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n614), .A2(new_n894), .A3(new_n623), .ZN(new_n895));
  NAND3_X1  g470(.A1(G299), .A2(new_n613), .A3(new_n608), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n614), .B2(new_n623), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n614), .A2(new_n623), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT101), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n896), .A4(new_n895), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n896), .A3(new_n895), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(KEYINPUT102), .A3(new_n893), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n847), .B(new_n631), .Z(new_n908));
  MUX2_X1   g483(.A(new_n907), .B(new_n905), .S(new_n908), .Z(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n909), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n715), .B(new_n601), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  XNOR2_X1  g491(.A(G305), .B(G166), .ZN(new_n917));
  MUX2_X1   g492(.A(new_n915), .B(new_n916), .S(new_n917), .Z(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n910), .B2(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n912), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n892), .B1(new_n920), .B2(new_n615), .ZN(G295));
  OAI21_X1  g496(.A(new_n892), .B1(new_n920), .B2(new_n615), .ZN(G331));
  XOR2_X1   g497(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n923));
  INV_X1    g498(.A(new_n905), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n579), .A2(new_n580), .A3(G301), .ZN(new_n925));
  NOR2_X1   g500(.A1(G171), .A2(G168), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n848), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT79), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n520), .B(new_n507), .C1(new_n508), .C2(new_n510), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n532), .A2(new_n527), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n539), .B1(new_n932), .B2(new_n537), .ZN(new_n933));
  AND4_X1   g508(.A1(new_n539), .A2(new_n537), .A3(new_n538), .A4(new_n524), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n536), .A2(KEYINPUT79), .A3(new_n540), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(G171), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G168), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G301), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n847), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n927), .A2(new_n928), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n847), .B1(new_n937), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT106), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n924), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n927), .A2(new_n940), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n944), .A2(KEYINPUT107), .B1(new_n907), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n937), .A2(new_n847), .A3(new_n939), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n947), .A2(new_n942), .A3(KEYINPUT106), .ZN(new_n948));
  INV_X1    g523(.A(new_n943), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n905), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n946), .A2(new_n918), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n887), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n918), .B1(new_n946), .B2(new_n952), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n927), .A2(new_n905), .A3(new_n940), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n941), .A2(new_n943), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n899), .A2(new_n903), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n917), .A2(new_n916), .ZN(new_n962));
  INV_X1    g537(.A(new_n917), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n915), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n953), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n923), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT107), .B(new_n905), .C1(new_n948), .C2(new_n949), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n945), .A2(new_n904), .A3(new_n906), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT107), .B1(new_n959), .B2(new_n905), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n970), .A2(new_n964), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n961), .A2(new_n964), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n887), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n976), .A2(new_n953), .A3(new_n957), .A4(new_n887), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT108), .B1(new_n967), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n977), .A3(KEYINPUT44), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n953), .A2(new_n957), .A3(new_n965), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n976), .A2(new_n887), .A3(new_n953), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(KEYINPUT43), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n980), .B(new_n981), .C1(new_n984), .C2(new_n923), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n497), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n464), .ZN(new_n991));
  INV_X1    g566(.A(new_n471), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n991), .B(G40), .C1(new_n992), .C2(new_n469), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n807), .B(G2067), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n771), .B(G1996), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n861), .A2(new_n731), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n728), .A2(new_n730), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n601), .B(new_n735), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G40), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n1002), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g579(.A(G2084), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n497), .A2(new_n987), .A3(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1003), .A2(new_n990), .A3(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(G168), .B(new_n1008), .C1(new_n1010), .C2(G1966), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n993), .B1(new_n989), .B2(new_n988), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1966), .B1(new_n1015), .B2(new_n1009), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1008), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n938), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT51), .A3(G8), .A4(new_n1011), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT123), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT62), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  OAI221_X1 g601(.A(G8), .B1(G288), .B2(new_n1026), .C1(new_n993), .C2(new_n988), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1031), .A3(KEYINPUT52), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1027), .B2(KEYINPUT52), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(G1981), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n593), .A2(new_n594), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n594), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n1038), .B2(new_n591), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT49), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n993), .B2(new_n988), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1025), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1034), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1032), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1042), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1046), .A2(new_n1052), .A3(KEYINPUT114), .A4(new_n1030), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n1056));
  OAI22_X1  g631(.A1(G166), .A2(new_n1055), .B1(KEYINPUT110), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n1058));
  NAND3_X1  g633(.A1(G303), .A2(G8), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT111), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(G2090), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1015), .A2(new_n1009), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n711), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1055), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1006), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n988), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n497), .A2(new_n1072), .A3(new_n987), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1003), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1068), .B1(G2090), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1060), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1064), .A2(new_n1069), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1015), .A2(new_n788), .A3(new_n1009), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1065), .A2(new_n795), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1080), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1079), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1010), .A2(KEYINPUT124), .A3(new_n788), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(KEYINPUT53), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1054), .A2(new_n1078), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT126), .B1(new_n1024), .B2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1054), .A2(new_n1078), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1014), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1022), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1094), .A2(new_n1098), .A3(new_n1099), .A4(new_n1091), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT62), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1093), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1043), .A2(G1976), .A3(G288), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1037), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1051), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1008), .B1(new_n1010), .B2(G1966), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1107), .A2(new_n581), .A3(G8), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1046), .A2(new_n1052), .A3(new_n1030), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT63), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1106), .B(new_n1111), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1108), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(KEYINPUT63), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1094), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1103), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1086), .A2(G301), .A3(new_n1090), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1084), .A2(new_n1085), .A3(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(KEYINPUT54), .C1(G301), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NOR4_X1   g697(.A1(new_n1084), .A2(new_n1085), .A3(G171), .A4(new_n1119), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1091), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1094), .A2(new_n1121), .A3(new_n1101), .A4(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n623), .B(KEYINPUT57), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT115), .B(G1956), .Z(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1074), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1015), .A2(new_n1009), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1126), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1126), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n993), .B1(new_n988), .B2(new_n1070), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1127), .B1(new_n1136), .B2(new_n1073), .ZN(new_n1137));
  AND4_X1   g712(.A1(new_n1003), .A2(new_n990), .A3(new_n1009), .A4(new_n1130), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1129), .A2(new_n1131), .A3(new_n1126), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT120), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1134), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n993), .A2(new_n988), .A3(KEYINPUT116), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT116), .B1(new_n993), .B2(new_n988), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT118), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1147), .A2(new_n1148), .A3(new_n1153), .A4(new_n1149), .ZN(new_n1154));
  INV_X1    g729(.A(G1996), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1010), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n561), .B(new_n1146), .C1(new_n1152), .C2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1139), .A2(KEYINPUT61), .A3(new_n1140), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1157), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n824), .B1(new_n1160), .B2(new_n1151), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1158), .B(new_n1159), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT122), .B1(new_n1145), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT121), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1134), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n809), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G1348), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1065), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1174), .A2(KEYINPUT117), .A3(new_n809), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1173), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1177), .A2(KEYINPUT60), .A3(new_n1181), .A4(new_n1179), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1183), .A2(new_n628), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1186), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1164), .A2(new_n1172), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1186), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1140), .A2(new_n628), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1132), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1125), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1001), .B1(new_n1117), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n995), .A2(new_n771), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n994), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n994), .A2(new_n1155), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT46), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT47), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1199), .B(KEYINPUT47), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(KEYINPUT127), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n807), .A2(new_n809), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n995), .A2(new_n996), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1206), .B1(new_n1207), .B2(new_n998), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n999), .A2(new_n994), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n994), .A2(new_n735), .A3(new_n601), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT48), .ZN(new_n1211));
  AOI22_X1  g786(.A1(new_n994), .A2(new_n1208), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1203), .A2(new_n1205), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1194), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g789(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n890), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1217), .A2(new_n984), .ZN(G308));
  OR2_X1    g792(.A1(new_n1217), .A2(new_n984), .ZN(G225));
endmodule


