//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975;
  AOI21_X1  g000(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT94), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G64gat), .Z(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT94), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n207), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n209), .A2(new_n203), .A3(new_n205), .A4(new_n204), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(G127gat), .ZN(new_n216));
  INV_X1    g015(.A(G22gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G15gat), .ZN(new_n218));
  INV_X1    g017(.A(G15gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT88), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n221), .A3(G1gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G8gat), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(new_n226), .A3(new_n231), .A4(new_n228), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT21), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n230), .B(new_n232), .C1(new_n211), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n216), .A2(new_n234), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G183gat), .B(G211gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n240), .B(new_n241), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OR3_X1    g042(.A1(new_n236), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n236), .B2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(KEYINPUT97), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(G99gat), .A3(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(G85gat), .ZN(new_n252));
  INV_X1    g051(.A(G92gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n249), .A2(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT7), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT96), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT96), .B1(new_n252), .B2(new_n253), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT96), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(G85gat), .A3(G92gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT7), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G99gat), .B(G106gat), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n254), .A2(new_n264), .A3(new_n256), .A4(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G50gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G43gat), .ZN(new_n269));
  INV_X1    g068(.A(G43gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G50gat), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT15), .ZN(new_n272));
  INV_X1    g071(.A(G36gat), .ZN(new_n273));
  INV_X1    g072(.A(G29gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT85), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G29gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n273), .A3(KEYINPUT14), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT14), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(G29gat), .B2(G36gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n272), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n272), .B(KEYINPUT86), .C1(new_n278), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT15), .B1(new_n269), .B2(new_n271), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n282), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT87), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT85), .B(G29gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n273), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT87), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n289), .A2(new_n290), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G232gat), .A2(G233gat), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n267), .A2(new_n296), .B1(KEYINPUT41), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299));
  INV_X1    g098(.A(new_n286), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n281), .B(new_n279), .C1(new_n292), .C2(new_n273), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT86), .B1(new_n301), .B2(new_n272), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n295), .B(new_n299), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n299), .B1(new_n287), .B2(new_n295), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n298), .B1(new_n306), .B2(new_n267), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT98), .ZN(new_n308));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n308), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n297), .A2(KEYINPUT41), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n312), .A2(new_n317), .A3(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n246), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n266), .A2(new_n211), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT99), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n263), .A2(new_n208), .A3(new_n210), .A4(new_n265), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n266), .A2(KEYINPUT99), .A3(new_n211), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT10), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT100), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n331));
  OR3_X1    g130(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n326), .B2(new_n331), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n323), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n323), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n336), .A3(new_n328), .ZN(new_n337));
  XNOR2_X1  g136(.A(G120gat), .B(G148gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT101), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT101), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n335), .A2(new_n343), .A3(new_n337), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n335), .A2(new_n337), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n322), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT93), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  INV_X1    g151(.A(G211gat), .ZN(new_n353));
  INV_X1    g152(.A(G218gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G211gat), .B(G218gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n360), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT26), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT27), .B(G183gat), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(KEYINPUT28), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  INV_X1    g168(.A(G183gat), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT27), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n374), .A2(KEYINPUT68), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT68), .B1(new_n374), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n368), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT69), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n365), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(KEYINPUT69), .B(new_n368), .C1(new_n376), .C2(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n370), .B2(new_n367), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n387));
  MUX2_X1   g186(.A(G183gat), .B(new_n387), .S(G190gat), .Z(new_n388));
  OAI211_X1 g187(.A(KEYINPUT65), .B(new_n383), .C1(new_n370), .C2(new_n367), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n362), .B1(new_n360), .B2(KEYINPUT23), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(KEYINPUT23), .B2(new_n360), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT25), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n362), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n399), .A2(KEYINPUT64), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n388), .A2(new_n384), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n399), .B2(KEYINPUT64), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n395), .A2(new_n396), .B1(new_n403), .B2(KEYINPUT25), .ZN(new_n404));
  INV_X1    g203(.A(G226gat), .ZN(new_n405));
  INV_X1    g204(.A(G233gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n382), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n406), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n382), .B2(new_n404), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n359), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n411), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n358), .A3(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(KEYINPUT37), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n420), .A2(new_n421), .B1(KEYINPUT37), .B2(new_n415), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT38), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n358), .A2(KEYINPUT82), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT37), .B1(new_n412), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n415), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(KEYINPUT82), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n423), .B(new_n419), .C1(new_n415), .C2(KEYINPUT37), .ZN(new_n428));
  OAI22_X1  g227(.A1(new_n422), .A2(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G162gat), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT2), .B1(new_n239), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G155gat), .B(G162gat), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G141gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(G148gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT74), .B(G141gat), .ZN(new_n439));
  INV_X1    g238(.A(G148gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G141gat), .B(G148gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(KEYINPUT2), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G113gat), .B(G120gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT1), .ZN(new_n447));
  XOR2_X1   g246(.A(G127gat), .B(G134gat), .Z(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(KEYINPUT4), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n444), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n447), .B(new_n448), .Z(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n445), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n442), .A2(new_n455), .A3(new_n444), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n450), .B(new_n454), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n449), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT76), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n452), .A2(new_n453), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n461), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT76), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n459), .A2(new_n472), .A3(new_n467), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G1gat), .B(G29gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT0), .ZN(new_n477));
  XNOR2_X1  g276(.A(G57gat), .B(G85gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n479), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n481), .A3(new_n474), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n473), .B1(new_n462), .B2(new_n470), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT78), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT6), .A4(new_n481), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n474), .A4(new_n481), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n412), .A2(new_n414), .A3(new_n418), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n484), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n429), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT3), .B1(new_n358), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n445), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n358), .B1(new_n457), .B2(new_n493), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT79), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(G228gat), .A3(G233gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(G228gat), .A2(G233gat), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT79), .B(new_n499), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n217), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT80), .ZN(new_n502));
  XOR2_X1   g301(.A(G78gat), .B(G106gat), .Z(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G50gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n498), .A2(new_n500), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G22gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n501), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n502), .A2(new_n508), .A3(new_n501), .A4(new_n505), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT39), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n459), .A2(new_n513), .A3(new_n467), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n514), .A2(new_n479), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n466), .A2(new_n468), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n461), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(KEYINPUT39), .C1(new_n460), .C2(new_n461), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n518), .A3(KEYINPUT40), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n519), .A2(new_n482), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT40), .B1(new_n515), .B2(new_n518), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT81), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT81), .ZN(new_n523));
  AOI211_X1 g322(.A(new_n523), .B(KEYINPUT40), .C1(new_n515), .C2(new_n518), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n420), .A2(KEYINPUT30), .A3(new_n490), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n415), .A2(KEYINPUT30), .A3(new_n419), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n512), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n489), .A2(new_n487), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n482), .A2(KEYINPUT77), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT77), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n485), .A2(new_n532), .A3(new_n481), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n531), .A2(new_n480), .A3(new_n533), .A4(new_n483), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n530), .A2(new_n534), .B1(new_n527), .B2(new_n526), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n492), .A2(new_n529), .B1(new_n535), .B2(new_n512), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n382), .A2(new_n449), .A3(new_n404), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n449), .B1(new_n382), .B2(new_n404), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G15gat), .B(G43gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G71gat), .B(G99gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT71), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n542), .A2(new_n550), .A3(KEYINPUT32), .A4(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n382), .A2(new_n404), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n453), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n382), .A2(new_n404), .A3(new_n449), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n538), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n553), .B1(new_n557), .B2(KEYINPUT33), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n545), .B1(new_n542), .B2(KEYINPUT32), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n542), .A2(KEYINPUT70), .A3(new_n546), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n538), .A3(new_n556), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n562), .A2(KEYINPUT72), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n562), .B2(KEYINPUT72), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n552), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n552), .B2(new_n561), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n537), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n561), .ZN(new_n571));
  INV_X1    g370(.A(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n561), .A3(new_n567), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT36), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n536), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n568), .A2(new_n569), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n512), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n573), .A2(new_n512), .A3(new_n579), .A4(new_n574), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n535), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n528), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n530), .B2(new_n484), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n512), .A3(new_n580), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n578), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n230), .A2(new_n232), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n296), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n230), .A2(KEYINPUT89), .A3(new_n232), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n592), .B(new_n593), .C1(new_n306), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT90), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT18), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n595), .B(new_n596), .C1(new_n304), .C2(new_n305), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n592), .A4(new_n593), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n601), .A2(KEYINPUT18), .A3(new_n592), .A4(new_n593), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n296), .B(new_n591), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n593), .B(KEYINPUT13), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n604), .B(new_n609), .C1(new_n611), .C2(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT92), .B1(new_n620), .B2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n350), .B1(new_n590), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n530), .A2(new_n534), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n528), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n573), .A2(new_n512), .A3(new_n574), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT83), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n630), .B2(new_n582), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n589), .B1(new_n631), .B2(new_n586), .ZN(new_n632));
  OAI221_X1 g431(.A(new_n576), .B1(new_n535), .B2(new_n512), .C1(new_n492), .C2(new_n529), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n625), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n349), .B1(new_n626), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n627), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT102), .B(G1gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1324gat));
  INV_X1    g440(.A(new_n528), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT16), .B(G8gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n231), .B1(new_n637), .B2(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT93), .B1(new_n634), .B2(new_n635), .ZN(new_n650));
  AOI211_X1 g449(.A(new_n350), .B(new_n625), .C1(new_n632), .C2(new_n633), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n642), .B(new_n348), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n643), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(KEYINPUT42), .ZN(new_n654));
  NOR4_X1   g453(.A1(new_n652), .A2(KEYINPUT103), .A3(new_n647), .A4(new_n643), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(G1325gat));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n219), .A3(new_n580), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n637), .A2(new_n577), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n659), .B2(new_n219), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n510), .A2(new_n511), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n637), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n246), .A2(new_n347), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n321), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n626), .B2(new_n636), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n669), .A2(KEYINPUT45), .A3(new_n638), .A4(new_n292), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n650), .B2(new_n651), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n638), .A2(new_n292), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n321), .B1(new_n632), .B2(new_n633), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n677), .B(new_n321), .C1(new_n632), .C2(new_n633), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n620), .A2(new_n622), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n679), .A2(new_n638), .A3(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n670), .B(new_n674), .C1(new_n683), .C2(new_n292), .ZN(G1328gat));
  NAND2_X1  g483(.A1(new_n642), .A2(new_n273), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n672), .A2(KEYINPUT46), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT46), .B1(new_n672), .B2(new_n685), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n679), .A2(new_n642), .A3(new_n682), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n686), .B(new_n687), .C1(new_n273), .C2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(new_n580), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n270), .B1(new_n672), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n576), .A2(new_n270), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n679), .A2(new_n682), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT47), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n691), .A2(new_n696), .A3(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1330gat));
  NAND3_X1  g497(.A1(new_n669), .A2(new_n268), .A3(new_n661), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n677), .B1(new_n590), .B2(new_n321), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n700), .A2(new_n701), .A3(new_n661), .A4(new_n682), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G50gat), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n699), .B2(new_n703), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(G1331gat));
  INV_X1    g506(.A(new_n347), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n322), .A2(new_n680), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n634), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n638), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n710), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n528), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  XNOR2_X1  g519(.A(new_n580), .B(KEYINPUT105), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(G71gat), .B1(new_n711), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n577), .A2(G71gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT50), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n711), .A2(G71gat), .A3(new_n577), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n715), .A2(new_n721), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(G71gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n661), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  INV_X1    g533(.A(new_n321), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n634), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n246), .A2(new_n680), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n737), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n708), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n252), .A3(new_n638), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n738), .A2(new_n708), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n679), .A2(new_n638), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n252), .B2(new_n744), .ZN(G1336gat));
  NAND4_X1  g544(.A1(new_n679), .A2(KEYINPUT106), .A3(new_n642), .A4(new_n743), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n700), .A2(new_n701), .A3(new_n642), .A4(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n749), .A3(G92gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n528), .A2(G92gat), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(new_n741), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n747), .A2(G92gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n740), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT51), .B1(new_n675), .B2(new_n737), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n347), .B(new_n751), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT52), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(G1337gat));
  NAND3_X1  g559(.A1(new_n679), .A2(new_n577), .A3(new_n743), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G99gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n741), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n690), .A2(G99gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(G1338gat));
  NAND4_X1  g564(.A1(new_n700), .A2(new_n701), .A3(new_n661), .A4(new_n743), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G106gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n512), .A2(G106gat), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n347), .B(new_n768), .C1(new_n755), .C2(new_n756), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT107), .B(KEYINPUT53), .Z(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n771), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1339gat));
  NOR3_X1   g574(.A1(new_n322), .A2(new_n680), .A3(new_n347), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n327), .A2(new_n328), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n331), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n779), .A2(new_n336), .A3(new_n332), .A4(new_n333), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n780), .A2(KEYINPUT54), .A3(new_n335), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n323), .C1(new_n329), .C2(new_n334), .ZN(new_n783));
  INV_X1    g582(.A(new_n340), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n777), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n780), .A2(new_n335), .A3(KEYINPUT54), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n784), .A4(new_n783), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n786), .A2(new_n345), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n604), .A2(new_n609), .A3(new_n621), .ZN(new_n790));
  INV_X1    g589(.A(new_n617), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n593), .B1(new_n601), .B2(new_n592), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n606), .A2(new_n607), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n735), .A2(new_n789), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n795), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n789), .A2(new_n680), .B1(new_n347), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(new_n735), .ZN(new_n801));
  INV_X1    g600(.A(new_n246), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n776), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n661), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n804), .A2(new_n638), .A3(new_n528), .A4(new_n580), .ZN(new_n805));
  INV_X1    g604(.A(G113gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n625), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n803), .A2(new_n627), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n581), .B2(new_n583), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n642), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n680), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n806), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n805), .A2(new_n813), .A3(new_n708), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n347), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n810), .A2(new_n817), .A3(new_n246), .ZN(new_n818));
  OAI21_X1  g617(.A(G127gat), .B1(new_n805), .B2(new_n802), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n642), .A2(new_n321), .ZN(new_n821));
  INV_X1    g620(.A(G134gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(KEYINPUT109), .B(KEYINPUT56), .Z(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n809), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n805), .B2(new_n321), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n809), .B2(new_n823), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT110), .ZN(G1343gat));
  AOI211_X1 g629(.A(new_n642), .B(new_n627), .C1(new_n570), .C2(new_n575), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n803), .B2(new_n512), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n512), .A2(new_n832), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n345), .A2(new_n788), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT111), .B1(new_n781), .B2(new_n785), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n787), .A2(new_n838), .A3(new_n784), .A4(new_n783), .ZN(new_n839));
  XOR2_X1   g638(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n836), .B(new_n841), .C1(new_n623), .C2(new_n624), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n347), .A2(new_n799), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n735), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n798), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n802), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n776), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n835), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n833), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n831), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n439), .B1(new_n852), .B2(new_n625), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n577), .A2(new_n512), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n808), .A2(new_n528), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n635), .A2(new_n436), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n853), .B(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n856), .A2(new_n857), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n680), .B(new_n831), .C1(new_n850), .C2(new_n851), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n439), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n859), .B2(new_n862), .ZN(G1344gat));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(G148gat), .C1(new_n852), .C2(new_n708), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n786), .A2(new_n345), .A3(new_n788), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n843), .B1(new_n681), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n321), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n246), .B1(new_n868), .B2(new_n798), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n834), .B1(new_n869), .B2(new_n776), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n348), .A2(new_n625), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n512), .B1(new_n846), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n347), .B1(new_n831), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n874), .B2(new_n831), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n440), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n864), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n877), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n865), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n856), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n440), .A3(new_n347), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1345gat));
  OAI21_X1  g684(.A(G155gat), .B1(new_n852), .B2(new_n802), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n883), .A2(new_n239), .A3(new_n246), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n852), .B2(new_n321), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n808), .A2(new_n430), .A3(new_n821), .A4(new_n855), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(KEYINPUT117), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n627), .A2(new_n642), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n721), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n804), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G169gat), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n625), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n801), .A2(new_n802), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n847), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n896), .B1(new_n630), .B2(new_n582), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n680), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n900), .A2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n904), .B2(new_n347), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT118), .ZN(new_n908));
  INV_X1    g707(.A(G176gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n898), .A2(new_n909), .A3(new_n708), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(G1349gat));
  AND2_X1   g710(.A1(new_n246), .A2(new_n366), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n902), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT119), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n902), .A2(new_n915), .A3(new_n903), .A4(new_n912), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n902), .A2(new_n512), .A3(new_n246), .A4(new_n897), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n914), .A2(new_n916), .B1(new_n917), .B2(G183gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT121), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT60), .B1(new_n918), .B2(KEYINPUT120), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n914), .A2(new_n916), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n917), .A2(G183gat), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n922), .A2(KEYINPUT120), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n918), .A2(KEYINPUT120), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT121), .A4(KEYINPUT60), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n925), .A2(new_n930), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n904), .A2(new_n367), .A3(new_n735), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT122), .Z(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n898), .B2(new_n321), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(G1351gat));
  NOR4_X1   g737(.A1(new_n803), .A2(new_n512), .A3(new_n577), .A4(new_n896), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n680), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n873), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n870), .B(KEYINPUT124), .C1(new_n872), .C2(KEYINPUT57), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n577), .A2(new_n896), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n944), .A2(new_n635), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G197gat), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n942), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NAND4_X1  g751(.A1(new_n944), .A2(new_n347), .A3(new_n945), .A4(new_n946), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n708), .A2(G204gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n954), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1353gat));
  NOR3_X1   g762(.A1(new_n577), .A2(new_n802), .A3(new_n896), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n353), .B1(new_n873), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT63), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n939), .A2(new_n353), .A3(new_n246), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1354gat));
  NAND4_X1  g767(.A1(new_n944), .A2(new_n735), .A3(new_n945), .A4(new_n946), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G218gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n939), .A2(new_n354), .A3(new_n735), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n974), .A3(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1355gat));
endmodule


