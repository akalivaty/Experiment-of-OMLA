//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n632, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT69), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G236), .A4(G238), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT71), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n468), .A3(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n462), .A2(new_n468), .A3(KEYINPUT72), .A4(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(G137), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n460), .A2(new_n461), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(G101), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  OAI221_X1 g063(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n477), .C2(G112), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT73), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n477), .A2(new_n481), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n481), .A2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(G124), .A2(new_n491), .B1(new_n492), .B2(G136), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n490), .A2(new_n493), .ZN(G162));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n481), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n475), .A2(new_n476), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n503), .A2(new_n462), .A3(new_n468), .A4(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G138), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n508), .B2(new_n481), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n501), .B1(new_n505), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n511), .A2(KEYINPUT74), .A3(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(G50), .A3(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(G75), .A2(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n518), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n517), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n517), .A2(new_n533), .A3(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n515), .A2(new_n516), .ZN(new_n538));
  INV_X1    g113(.A(new_n512), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n538), .A2(new_n539), .A3(new_n527), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G89), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n544));
  AND2_X1   g119(.A1(G63), .A2(G651), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n527), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT76), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n536), .ZN(new_n549));
  OAI21_X1  g124(.A(G51), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n550), .A2(new_n551), .A3(new_n541), .A4(new_n546), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G168));
  AOI22_X1  g128(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n554), .A2(new_n555), .A3(new_n514), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n554), .B2(new_n514), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(new_n557), .B1(G90), .B2(new_n540), .ZN(new_n558));
  OAI21_X1  g133(.A(G52), .B1(new_n549), .B2(new_n534), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(new_n540), .A2(G81), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n514), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n563), .A2(new_n566), .A3(new_n514), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n562), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n549), .A2(new_n534), .ZN(new_n569));
  INV_X1    g144(.A(G43), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(G188));
  NAND3_X1  g152(.A1(new_n538), .A2(G543), .A3(new_n539), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n517), .A2(new_n581), .A3(G53), .A4(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n517), .A2(G91), .A3(new_n527), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n522), .B2(new_n523), .ZN(new_n586));
  AND2_X1   g161(.A1(G78), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n583), .A2(new_n589), .ZN(G299));
  INV_X1    g165(.A(G168), .ZN(G286));
  OAI21_X1  g166(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n592));
  INV_X1    g167(.A(G49), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n592), .B1(new_n578), .B2(new_n593), .C1(new_n594), .C2(new_n528), .ZN(G288));
  AND2_X1   g170(.A1(G48), .A2(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n538), .A2(new_n539), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n517), .A2(KEYINPUT79), .A3(new_n596), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n599), .A2(new_n600), .B1(new_n540), .B2(G86), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n514), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(G305));
  OAI21_X1  g180(.A(G47), .B1(new_n549), .B2(new_n534), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n522), .A2(new_n523), .ZN(new_n608));
  INV_X1    g183(.A(G60), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(G85), .A2(new_n540), .B1(new_n610), .B2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n606), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n528), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n608), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n616), .A2(new_n619), .B1(G651), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(G54), .B1(new_n549), .B2(new_n534), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n614), .B1(new_n615), .B2(new_n627), .ZN(G284));
  AOI21_X1  g203(.A(new_n614), .B1(new_n615), .B2(new_n627), .ZN(G321));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  MUX2_X1   g208(.A(new_n630), .B(new_n632), .S(new_n633), .Z(G297));
  MUX2_X1   g209(.A(new_n630), .B(new_n632), .S(new_n633), .Z(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n626), .B1(new_n636), .B2(G860), .ZN(G148));
  OAI21_X1  g212(.A(KEYINPUT82), .B1(new_n572), .B2(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n626), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  MUX2_X1   g215(.A(KEYINPUT82), .B(new_n638), .S(new_n640), .Z(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g217(.A1(new_n462), .A2(new_n468), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(new_n485), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AOI22_X1  g224(.A1(G123), .A2(new_n491), .B1(new_n492), .B2(G135), .ZN(new_n650));
  OAI221_X1 g225(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n477), .C2(G111), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(G156));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n658), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n672), .B(new_n678), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n674), .C1(new_n671), .C2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n671), .A3(new_n673), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n686), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n686), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  NOR2_X1   g278(.A1(G29), .A2(G35), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G162), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT29), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G2090), .Z(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(G171), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G5), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n713));
  INV_X1    g288(.A(G1348), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n626), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G4), .B2(G16), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n708), .A2(G19), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n572), .B2(new_n708), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1341), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n707), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  OAI22_X1  g296(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n708), .A2(G20), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT23), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G299), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(G160), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n726), .B1(G2084), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n721), .A2(new_n722), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT25), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n643), .A2(G127), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n477), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n737), .B(new_n740), .C1(G139), .C2(new_n492), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n731), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2072), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n731), .A2(G26), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT28), .Z(new_n745));
  AOI22_X1  g320(.A1(G128), .A2(new_n491), .B1(new_n492), .B2(G140), .ZN(new_n746));
  OAI221_X1 g321(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n477), .C2(G116), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n751), .A2(new_n731), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n652), .B2(new_n731), .ZN(new_n755));
  NAND2_X1  g330(.A1(G164), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G27), .B2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT93), .B(G2078), .Z(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n750), .B(new_n759), .C1(new_n757), .C2(new_n758), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n743), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n710), .A2(new_n711), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n708), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n708), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n761), .B(new_n762), .C1(G1966), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G1966), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n491), .A2(G129), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n492), .A2(G141), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n485), .A2(new_n772), .A3(G105), .ZN(new_n773));
  INV_X1    g348(.A(G105), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT87), .B1(new_n484), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n770), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n770), .B2(new_n777), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT89), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G29), .B2(G32), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT90), .B2(new_n783), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT91), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n732), .A2(G2084), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT86), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n734), .A2(new_n766), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G23), .B(G288), .S(G16), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT33), .B(G1976), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n708), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n708), .ZN(new_n798));
  INV_X1    g373(.A(G1971), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT32), .B(G1981), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT85), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n731), .A2(G25), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n491), .A2(G119), .ZN(new_n812));
  OAI221_X1 g387(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n477), .C2(G107), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n492), .A2(G131), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n811), .B1(new_n816), .B2(new_n731), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G290), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n708), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n708), .B2(G24), .ZN(new_n822));
  INV_X1    g397(.A(G1986), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n809), .A2(new_n810), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n793), .B1(new_n827), .B2(new_n828), .ZN(G311));
  XNOR2_X1  g404(.A(new_n826), .B(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(new_n793), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(G150));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n608), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n514), .B1(new_n835), .B2(KEYINPUT94), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(new_n833), .C1(new_n608), .C2(new_n834), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n836), .A2(new_n838), .B1(G93), .B2(new_n540), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n840));
  OAI21_X1  g415(.A(G55), .B1(new_n549), .B2(new_n534), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n842), .A2(new_n843), .B1(new_n571), .B2(new_n568), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n572), .A2(new_n841), .A3(new_n839), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n626), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n741), .A2(new_n781), .ZN(new_n857));
  INV_X1    g432(.A(new_n782), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n741), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n748), .B(G164), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n491), .A2(G130), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT96), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n492), .A2(G142), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n477), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n861), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n645), .B(new_n815), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n860), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G160), .B(G162), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n652), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n859), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n875), .B1(new_n873), .B2(new_n876), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n856), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n882), .A2(KEYINPUT97), .A3(new_n878), .A4(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g460(.A(new_n846), .B(new_n639), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n625), .A2(G299), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n631), .A2(new_n624), .A3(new_n623), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(KEYINPUT98), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n891), .A2(KEYINPUT98), .ZN(new_n897));
  XNOR2_X1  g472(.A(G290), .B(G305), .ZN(new_n898));
  XNOR2_X1  g473(.A(G288), .B(G303), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT42), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n896), .B2(new_n897), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n842), .A2(new_n843), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n905), .ZN(G295));
  OAI21_X1  g481(.A(new_n904), .B1(G868), .B2(new_n905), .ZN(G331));
  NAND2_X1  g482(.A1(new_n839), .A2(new_n841), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT95), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n572), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n908), .A2(new_n571), .A3(new_n568), .ZN(new_n912));
  NAND3_X1  g487(.A1(G301), .A2(new_n548), .A3(new_n552), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G301), .B1(new_n552), .B2(new_n548), .ZN(new_n915));
  OAI22_X1  g490(.A1(new_n911), .A2(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(G171), .A2(G168), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n844), .A2(new_n917), .A3(new_n845), .A4(new_n913), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n916), .A2(new_n918), .A3(new_n890), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n916), .A2(new_n918), .B1(new_n893), .B2(new_n894), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n921), .B2(new_n900), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(new_n918), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n893), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT101), .A4(new_n892), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n894), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n924), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(new_n919), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n922), .B(new_n923), .C1(new_n932), .C2(new_n900), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  INV_X1    g509(.A(new_n900), .ZN(new_n935));
  INV_X1    g510(.A(new_n919), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n924), .A2(new_n929), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n925), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n938), .B2(new_n930), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n922), .A4(new_n923), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n922), .B1(new_n900), .B2(new_n921), .ZN(new_n942));
  INV_X1    g517(.A(new_n923), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n934), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n922), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n949), .B(KEYINPUT44), .C1(new_n942), .C2(new_n943), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n465), .A2(new_n467), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n477), .A3(G138), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n643), .A2(new_n953), .B1(new_n955), .B2(KEYINPUT4), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n956), .B2(new_n501), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT45), .B1(new_n957), .B2(KEYINPUT104), .ZN(new_n958));
  INV_X1    g533(.A(G101), .ZN(new_n959));
  OAI221_X1 g534(.A(G40), .B1(new_n959), .B2(new_n484), .C1(new_n480), .C2(new_n481), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n474), .B2(new_n478), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n958), .B(new_n961), .C1(KEYINPUT104), .C2(new_n957), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n820), .A2(new_n823), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT106), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n820), .A2(new_n823), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT107), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n858), .A2(G1996), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n748), .A2(G2067), .ZN(new_n974));
  INV_X1    g549(.A(G2067), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n746), .A2(new_n975), .A3(new_n747), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n781), .B2(G1996), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n816), .A2(new_n818), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n816), .A2(new_n818), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n973), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n972), .B1(new_n967), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n952), .C1(new_n956), .C2(new_n501), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n961), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n711), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT122), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n952), .C1(new_n956), .C2(new_n501), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(G164), .B2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G2078), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n961), .A2(new_n989), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n987), .A2(new_n988), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n988), .B1(new_n987), .B2(new_n994), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n961), .A2(new_n989), .A3(new_n991), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT108), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n961), .A2(new_n989), .A3(new_n991), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G2078), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n995), .A2(new_n996), .B1(new_n1001), .B2(KEYINPUT53), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G171), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT123), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n958), .B1(KEYINPUT104), .B2(new_n957), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n989), .A2(G40), .A3(new_n993), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n487), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1007), .A2(new_n1009), .B1(new_n711), .B2(new_n986), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1001), .B2(KEYINPUT53), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(G171), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1006), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(KEYINPUT125), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT125), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1010), .B(new_n1016), .C1(KEYINPUT53), .C2(new_n1001), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G171), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1002), .A2(G171), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1013), .A2(new_n1014), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G286), .A2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n961), .A2(new_n989), .A3(new_n991), .ZN(new_n1026));
  INV_X1    g601(.A(G2084), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n961), .A2(new_n984), .A3(new_n985), .A4(new_n1027), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1026), .A2(G1966), .B1(new_n1028), .B2(KEYINPUT115), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1025), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n997), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1024), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1036), .A3(G168), .ZN(new_n1038));
  AND2_X1   g613(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1037), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  INV_X1    g620(.A(G1956), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n986), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n583), .A2(KEYINPUT116), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n1049));
  NAND3_X1  g624(.A1(G299), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n583), .B(new_n589), .C1(KEYINPUT116), .C2(KEYINPUT57), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT56), .B(G2072), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n961), .A2(new_n989), .A3(new_n991), .A4(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1047), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1045), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT118), .B(new_n1045), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1052), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1047), .A2(KEYINPUT117), .A3(new_n1054), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1055), .A2(new_n1045), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n997), .A2(G1996), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n505), .A2(new_n509), .ZN(new_n1070));
  INV_X1    g645(.A(new_n501), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1384), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1069), .B1(new_n961), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n572), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT59), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(new_n572), .C1(new_n1068), .C2(new_n1073), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1066), .A2(new_n1067), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n986), .A2(new_n714), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n961), .A2(new_n975), .A3(new_n1072), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT60), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT119), .B1(new_n1081), .B2(new_n625), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  INV_X1    g658(.A(new_n960), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n479), .A2(new_n1084), .A3(new_n1072), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1086), .A2(new_n975), .B1(new_n986), .B2(new_n714), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(new_n626), .C1(new_n1087), .C2(KEYINPUT60), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1082), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(KEYINPUT60), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1061), .A2(new_n1078), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1055), .A2(new_n625), .A3(new_n1087), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1044), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1976), .ZN(new_n1098));
  OR2_X1    g673(.A1(G288), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G8), .ZN(new_n1100));
  AOI211_X1 g675(.A(KEYINPUT111), .B(new_n1100), .C1(new_n961), .C2(new_n1072), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1085), .B2(G8), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n1106));
  INV_X1    g681(.A(G1981), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n517), .A2(G86), .A3(new_n527), .ZN(new_n1108));
  AND4_X1   g683(.A1(KEYINPUT79), .A2(new_n538), .A3(new_n539), .A4(new_n596), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT79), .B1(new_n517), .B2(new_n596), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n603), .B1(new_n1111), .B2(KEYINPUT113), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1107), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT112), .B(G1981), .Z(new_n1116));
  NOR2_X1   g691(.A1(G305), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1106), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n604), .B1(new_n601), .B2(new_n1113), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1114), .ZN(new_n1120));
  OAI21_X1  g695(.A(G1981), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(G305), .A2(new_n1116), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT49), .A3(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1118), .B(new_n1123), .C1(new_n1101), .C2(new_n1103), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT52), .B1(G288), .B2(new_n1098), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1099), .B(new_n1125), .C1(new_n1101), .C2(new_n1103), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1105), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(G303), .A2(G8), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT55), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT110), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(KEYINPUT110), .A3(new_n1129), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT109), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT109), .ZN(new_n1135));
  NAND4_X1  g710(.A1(G303), .A2(new_n1135), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n998), .A2(new_n799), .A3(new_n1000), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n986), .A2(G2090), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1100), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1127), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(KEYINPUT114), .A3(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G8), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT114), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1137), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1141), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1142), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1023), .A2(new_n1097), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1140), .ZN(new_n1151));
  NOR2_X1   g726(.A1(G288), .A2(G1976), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1117), .B1(new_n1124), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1151), .A2(new_n1127), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1041), .A2(G286), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1141), .A2(new_n1146), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1137), .B1(new_n1160), .B2(new_n1100), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1141), .A2(new_n1156), .A3(KEYINPUT63), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1155), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1150), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(new_n1044), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1038), .A2(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1167), .B(KEYINPUT62), .C1(new_n1168), .C2(new_n1037), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1044), .A2(new_n1165), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT124), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1141), .A2(new_n1146), .A3(new_n1142), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n982), .B1(new_n1164), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n973), .A2(new_n978), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n976), .B1(new_n1179), .B2(new_n980), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n967), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n981), .A2(new_n967), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n967), .A2(new_n969), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT48), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1181), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n966), .A2(G1996), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT46), .Z(new_n1190));
  OAI21_X1  g765(.A(new_n967), .B1(new_n781), .B2(new_n977), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1192), .A2(KEYINPUT47), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(KEYINPUT47), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1178), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g771(.A1(G227), .A2(new_n458), .ZN(new_n1198));
  XOR2_X1   g772(.A(new_n1198), .B(KEYINPUT127), .Z(new_n1199));
  NOR3_X1   g773(.A1(G229), .A2(G401), .A3(new_n1199), .ZN(new_n1200));
  AND3_X1   g774(.A1(new_n945), .A2(new_n884), .A3(new_n1200), .ZN(G308));
  NAND3_X1  g775(.A1(new_n945), .A2(new_n884), .A3(new_n1200), .ZN(G225));
endmodule


