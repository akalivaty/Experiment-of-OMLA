//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  OR3_X1    g001(.A1(new_n202), .A2(G29gat), .A3(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT87), .B(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  AOI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n207), .A2(new_n209), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n214), .A2(KEYINPUT17), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(new_n220), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n214), .A2(KEYINPUT17), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT90), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n214), .B(new_n220), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n226), .B(KEYINPUT13), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G197gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT11), .B(G169gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  XOR2_X1   g040(.A(new_n229), .B(KEYINPUT91), .Z(new_n242));
  NOR2_X1   g041(.A1(new_n235), .A2(new_n241), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n236), .A2(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G85gat), .ZN(new_n245));
  INV_X1    g044(.A(G92gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT96), .ZN(new_n247));
  AOI211_X1 g046(.A(new_n245), .B(new_n246), .C1(new_n247), .C2(KEYINPUT7), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n247), .B2(KEYINPUT7), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT7), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT96), .B(new_n250), .C1(new_n245), .C2(new_n246), .ZN(new_n251));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252));
  AOI22_X1  g051(.A1(KEYINPUT8), .A2(new_n252), .B1(new_n245), .B2(new_n246), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G99gat), .B(G106gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n224), .A2(new_n222), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT41), .ZN(new_n258));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259));
  OAI221_X1 g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .C1(new_n214), .C2(new_n256), .ZN(new_n260));
  XNOR2_X1  g059(.A(G190gat), .B(G218gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n258), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT97), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(KEYINPUT97), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n262), .B1(new_n269), .B2(new_n267), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G57gat), .B(G64gat), .Z(new_n272));
  INV_X1    g071(.A(KEYINPUT9), .ZN(new_n273));
  INV_X1    g072(.A(G71gat), .ZN(new_n274));
  INV_X1    g073(.A(G78gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(KEYINPUT92), .A3(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G71gat), .B(G78gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n281), .B(KEYINPUT93), .Z(new_n282));
  XOR2_X1   g081(.A(G127gat), .B(G155gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT20), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n282), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G211gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT95), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n279), .B(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n220), .B1(new_n289), .B2(new_n280), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n291));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n290), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n287), .B(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n271), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n255), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT98), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n254), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n299), .B2(new_n254), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT99), .ZN(new_n302));
  INV_X1    g101(.A(new_n279), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n254), .A2(new_n255), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(KEYINPUT99), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n256), .A2(new_n279), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n308));
  AND3_X1   g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n289), .A2(new_n310), .A3(new_n256), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT101), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n297), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n306), .A2(new_n307), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n297), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G120gat), .B(G148gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT102), .ZN(new_n318));
  XOR2_X1   g117(.A(G176gat), .B(G204gat), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n320), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n327), .A2(new_n328), .B1(new_n329), .B2(KEYINPUT28), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n329), .B2(KEYINPUT28), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n327), .A2(KEYINPUT69), .A3(new_n333), .A4(new_n328), .ZN(new_n334));
  AND2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  INV_X1    g134(.A(G169gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n335), .B1(new_n338), .B2(KEYINPUT26), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(KEYINPUT26), .B2(new_n338), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n344), .A2(G169gat), .A3(G176gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n345), .B2(new_n335), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n332), .ZN(new_n348));
  NAND3_X1  g147(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT67), .B(new_n351), .C1(new_n338), .C2(new_n344), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n338), .B2(new_n344), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n346), .A2(new_n350), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n348), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT65), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n358), .A2(new_n359), .B1(new_n332), .B2(new_n347), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n335), .B1(new_n338), .B2(new_n344), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n344), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n336), .ZN(new_n369));
  NAND2_X1  g168(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n362), .A2(new_n365), .A3(new_n373), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n342), .B(new_n356), .C1(new_n374), .C2(new_n353), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n371), .B(new_n366), .C1(new_n363), .C2(new_n364), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT65), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n353), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT68), .B1(new_n378), .B2(new_n355), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n341), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G113gat), .ZN(new_n381));
  INV_X1    g180(.A(G120gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT1), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n381), .B2(new_n382), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n385), .A2(KEYINPUT70), .B1(G127gat), .B2(G134gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(G127gat), .B2(G134gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n384), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n372), .B1(KEYINPUT65), .B2(new_n361), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT25), .B1(new_n391), .B2(new_n365), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n342), .B1(new_n392), .B2(new_n356), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT68), .A3(new_n355), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n388), .A3(new_n341), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G227gat), .ZN(new_n398));
  INV_X1    g197(.A(G233gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT71), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT71), .ZN(new_n402));
  INV_X1    g201(.A(new_n400), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n402), .B(new_n403), .C1(new_n390), .C2(new_n396), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n326), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G15gat), .B(G43gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n388), .B1(new_n395), .B2(new_n341), .ZN(new_n411));
  INV_X1    g210(.A(new_n341), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n389), .B(new_n412), .C1(new_n393), .C2(new_n394), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n400), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n402), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n397), .A2(KEYINPUT71), .A3(new_n400), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n410), .B1(new_n417), .B2(KEYINPUT32), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT72), .A3(new_n326), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n407), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n417), .B(KEYINPUT32), .C1(new_n326), .C2(new_n410), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n420), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n397), .A2(new_n400), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT32), .B1(new_n401), .B2(new_n404), .ZN(new_n428));
  INV_X1    g227(.A(new_n410), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT33), .B1(new_n415), .B2(new_n416), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n428), .B(new_n429), .C1(new_n430), .C2(KEYINPUT72), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n405), .A2(new_n406), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n422), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n425), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT73), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n426), .B1(new_n423), .B2(new_n424), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n425), .A3(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT73), .A3(KEYINPUT36), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT81), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT31), .ZN(new_n446));
  INV_X1    g245(.A(G50gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n450));
  OR2_X1    g249(.A1(G197gat), .A2(G204gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(G197gat), .A2(G204gat), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT74), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n453), .A2(new_n454), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n456), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT75), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT79), .B(G148gat), .Z(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G141gat), .ZN(new_n464));
  INV_X1    g263(.A(G148gat), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n465), .A2(G141gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(G155gat), .A2(G162gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(KEYINPUT2), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n468), .ZN(new_n474));
  AND2_X1   g273(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n475));
  NOR2_X1   g274(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT78), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n465), .A2(G141gat), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n477), .A2(new_n478), .B1(new_n466), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n474), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n462), .B1(new_n486), .B2(KEYINPUT29), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n449), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT29), .B1(new_n457), .B2(new_n459), .ZN(new_n490));
  OAI22_X1  g289(.A1(new_n490), .A2(KEYINPUT3), .B1(new_n473), .B2(new_n482), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n487), .B(new_n491), .C1(new_n488), .C2(new_n449), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(G22gat), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n448), .B1(new_n496), .B2(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n494), .ZN(new_n498));
  INV_X1    g297(.A(G22gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n500), .A2(KEYINPUT83), .A3(new_n495), .A4(new_n448), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n388), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n483), .A2(new_n388), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(KEYINPUT80), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT5), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT3), .B1(new_n473), .B2(new_n482), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n485), .A2(new_n513), .A3(new_n389), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n505), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n511), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(KEYINPUT5), .A3(new_n511), .A4(new_n514), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G1gat), .B(G29gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT0), .ZN(new_n524));
  XNOR2_X1  g323(.A(G57gat), .B(G85gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528));
  INV_X1    g327(.A(new_n526), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n519), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n530), .A2(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(G226gat), .A2(G233gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT29), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n412), .B1(new_n378), .B2(new_n355), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n380), .A2(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n462), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n378), .A2(new_n355), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n341), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n535), .ZN(new_n541));
  NAND2_X1  g340(.A1(G226gat), .A2(G233gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n380), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n462), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G8gat), .B(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT76), .ZN(new_n548));
  XNOR2_X1  g347(.A(G64gat), .B(G92gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  NOR2_X1   g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n553), .B1(new_n546), .B2(new_n550), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n504), .A2(new_n533), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n550), .B1(new_n546), .B2(KEYINPUT37), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n538), .B2(new_n545), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT85), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n561), .B1(new_n537), .B2(new_n544), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n462), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n565), .A2(new_n566), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT38), .B1(new_n569), .B2(new_n564), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n563), .A2(KEYINPUT38), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n530), .A2(new_n528), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n529), .B1(new_n519), .B2(new_n521), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT84), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT84), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n527), .A2(new_n575), .A3(new_n528), .A4(new_n530), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n532), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n551), .ZN(new_n578));
  INV_X1    g377(.A(new_n557), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n520), .A2(new_n514), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n510), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n508), .A2(new_n511), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT39), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n584), .A3(new_n510), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n526), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT40), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n530), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n587), .B2(new_n586), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n571), .A2(new_n578), .B1(new_n579), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n559), .B1(new_n590), .B2(new_n504), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n439), .A2(new_n443), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n427), .A2(new_n436), .ZN(new_n593));
  INV_X1    g392(.A(new_n504), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT86), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n557), .A2(new_n577), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n557), .B2(new_n577), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT35), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n533), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n579), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n440), .A2(new_n441), .A3(new_n601), .A4(new_n594), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT35), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n244), .B(new_n325), .C1(new_n592), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n600), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT103), .B(G1gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(G1324gat));
  AND2_X1   g407(.A1(new_n605), .A2(new_n579), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n219), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT104), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT16), .B(G8gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT42), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(G1325gat));
  INV_X1    g414(.A(G15gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n616), .A3(new_n593), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT36), .B1(new_n442), .B2(KEYINPUT73), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n619));
  AOI211_X1 g418(.A(new_n619), .B(new_n438), .C1(new_n440), .C2(new_n441), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n605), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n623), .B2(new_n616), .ZN(G1326gat));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n504), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT43), .B(G22gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(G1327gat));
  AND2_X1   g426(.A1(new_n268), .A2(new_n270), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(new_n592), .B2(new_n604), .ZN(new_n629));
  INV_X1    g428(.A(new_n295), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n244), .A2(new_n630), .A3(new_n323), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n600), .A3(new_n205), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT45), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT105), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n592), .A2(new_n636), .A3(new_n604), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n592), .B2(new_n604), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n271), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n629), .A2(new_n639), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n631), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(KEYINPUT106), .B(new_n631), .C1(new_n641), .C2(new_n642), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n646), .A2(new_n648), .A3(new_n533), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n635), .B1(new_n649), .B2(new_n205), .ZN(G1328gat));
  NOR3_X1   g449(.A1(new_n632), .A2(G36gat), .A3(new_n557), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT46), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n646), .A2(new_n648), .A3(new_n557), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n206), .ZN(G1329gat));
  OAI21_X1  g453(.A(G43gat), .B1(new_n643), .B2(new_n621), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n632), .A2(G43gat), .A3(new_n442), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT47), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n645), .A2(new_n622), .A3(new_n647), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n660), .B2(G43gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n661), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g461(.A(G50gat), .B1(new_n643), .B2(new_n594), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n633), .A2(KEYINPUT107), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n447), .B(new_n504), .C1(new_n632), .C2(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n663), .B(KEYINPUT48), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n645), .A2(new_n504), .A3(new_n647), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(G50gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n670), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g470(.A1(new_n637), .A2(new_n638), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n244), .A2(new_n296), .A3(new_n323), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n533), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT108), .B(G57gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1332gat));
  AND2_X1   g476(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n557), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT109), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1333gat));
  NAND3_X1  g485(.A1(new_n678), .A2(new_n274), .A3(new_n593), .ZN(new_n687));
  OAI21_X1  g486(.A(G71gat), .B1(new_n674), .B2(new_n621), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n594), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n275), .ZN(G1335gat));
  NAND2_X1  g491(.A1(new_n244), .A2(new_n295), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n578), .A2(new_n571), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n579), .A2(new_n589), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n558), .B1(new_n697), .B2(new_n594), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n618), .A2(new_n620), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n442), .A2(new_n504), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n700), .A2(new_n598), .B1(new_n602), .B2(KEYINPUT35), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n271), .B(new_n694), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n629), .A2(KEYINPUT51), .A3(new_n694), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n706), .A2(new_n245), .A3(new_n600), .A4(new_n323), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n693), .A2(new_n324), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n641), .ZN(new_n710));
  INV_X1    g509(.A(new_n642), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n600), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n713), .B2(new_n245), .ZN(G1336gat));
  INV_X1    g513(.A(new_n706), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n323), .A2(new_n579), .A3(new_n246), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n712), .A2(new_n579), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n246), .ZN(new_n721));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n246), .B1(new_n712), .B2(new_n579), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(G1337gat));
  AND2_X1   g524(.A1(new_n712), .A2(new_n622), .ZN(new_n726));
  INV_X1    g525(.A(G99gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n593), .A2(new_n727), .A3(new_n323), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n726), .A2(new_n727), .B1(new_n715), .B2(new_n728), .ZN(G1338gat));
  OAI211_X1 g528(.A(new_n504), .B(new_n708), .C1(new_n641), .C2(new_n642), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G106gat), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n324), .A2(new_n594), .A3(G106gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n706), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT53), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n592), .A2(new_n604), .ZN(new_n736));
  AND4_X1   g535(.A1(KEYINPUT51), .A2(new_n736), .A3(new_n271), .A4(new_n694), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT51), .B1(new_n629), .B2(new_n694), .ZN(new_n738));
  OAI211_X1 g537(.A(KEYINPUT111), .B(new_n732), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT111), .B1(new_n706), .B2(new_n732), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT112), .B1(new_n743), .B2(new_n731), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n732), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n704), .B2(new_n705), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT53), .B1(new_n748), .B2(KEYINPUT111), .ZN(new_n749));
  AND4_X1   g548(.A1(KEYINPUT112), .A2(new_n731), .A3(new_n746), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(G1339gat));
  NAND2_X1  g550(.A1(new_n242), .A2(new_n243), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n230), .A2(new_n235), .ZN(new_n753));
  INV_X1    g552(.A(new_n241), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n325), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n311), .B(KEYINPUT101), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n759), .A3(G230gat), .A4(G233gat), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n314), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n320), .B1(new_n314), .B2(KEYINPUT54), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n314), .A2(KEYINPUT54), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n314), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n764), .A2(KEYINPUT55), .A3(new_n320), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n766), .A3(new_n321), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n225), .A2(new_n226), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n232), .A2(new_n233), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n240), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n770), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n244), .A2(new_n767), .B1(new_n324), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n628), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n763), .A2(new_n321), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n271), .A3(new_n766), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n775), .A2(new_n771), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n756), .B1(new_n777), .B2(new_n295), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n533), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n700), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n557), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n244), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n381), .ZN(G1340gat));
  NOR2_X1   g582(.A1(new_n781), .A2(new_n324), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(new_n382), .ZN(G1341gat));
  NOR2_X1   g584(.A1(new_n781), .A2(new_n295), .ZN(new_n786));
  INV_X1    g585(.A(G127gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT113), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n786), .B(new_n788), .Z(G1342gat));
  INV_X1    g588(.A(G134gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n271), .A2(new_n557), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT114), .Z(new_n792));
  NAND3_X1  g591(.A1(new_n780), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT56), .Z(new_n794));
  OAI21_X1  g593(.A(G134gat), .B1(new_n781), .B2(new_n628), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1343gat));
  AND2_X1   g595(.A1(new_n779), .A2(KEYINPUT115), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n504), .B1(new_n779), .B2(KEYINPUT115), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(new_n798), .A3(new_n622), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n244), .A2(G141gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n557), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n579), .A2(new_n533), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n755), .A2(new_n766), .A3(new_n774), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n752), .A2(new_n770), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n323), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n271), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n775), .A2(new_n771), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n295), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n756), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n594), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(KEYINPUT57), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812));
  AOI211_X1 g611(.A(new_n812), .B(new_n594), .C1(new_n808), .C2(new_n809), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n621), .B(new_n802), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G141gat), .B1(new_n814), .B2(new_n244), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n801), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT58), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n818), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1344gat));
  AND2_X1   g619(.A1(new_n799), .A2(new_n557), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n463), .A3(new_n323), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n463), .A2(KEYINPUT59), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n814), .B2(new_n324), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n628), .A2(new_n767), .A3(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n775), .A2(KEYINPUT117), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n804), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n630), .B1(new_n830), .B2(new_n773), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n504), .B1(new_n831), .B2(new_n756), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n813), .B1(new_n812), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n621), .A2(new_n323), .A3(new_n802), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(KEYINPUT118), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n465), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT118), .B1(new_n833), .B2(new_n834), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n827), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n822), .B1(new_n826), .B2(new_n838), .ZN(G1345gat));
  INV_X1    g638(.A(G155gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n840), .A3(new_n630), .ZN(new_n841));
  OAI21_X1  g640(.A(G155gat), .B1(new_n814), .B2(new_n295), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1346gat));
  INV_X1    g642(.A(G162gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n799), .A2(new_n844), .A3(new_n792), .ZN(new_n845));
  OAI21_X1  g644(.A(G162gat), .B1(new_n814), .B2(new_n628), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1347gat));
  INV_X1    g646(.A(new_n778), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n557), .A2(new_n600), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n700), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n244), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(G169gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n369), .A2(new_n370), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1348gat));
  NOR2_X1   g653(.A1(new_n850), .A2(new_n324), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(new_n337), .ZN(G1349gat));
  OR2_X1    g655(.A1(new_n850), .A2(new_n295), .ZN(new_n857));
  INV_X1    g656(.A(G183gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n327), .B2(new_n857), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1350gat));
  NOR2_X1   g661(.A1(new_n850), .A2(new_n628), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n328), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT61), .Z(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n328), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT119), .Z(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1351gat));
  NAND2_X1  g667(.A1(new_n621), .A2(new_n849), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n778), .A2(new_n869), .A3(new_n594), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n244), .A2(G197gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  MUX2_X1   g674(.A(new_n810), .B(new_n832), .S(new_n812), .Z(new_n876));
  OR2_X1    g675(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G197gat), .B1(new_n879), .B2(new_n244), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT122), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n875), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1352gat));
  XOR2_X1   g684(.A(KEYINPUT123), .B(G204gat), .Z(new_n886));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n323), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT62), .Z(new_n888));
  NOR2_X1   g687(.A1(new_n879), .A2(new_n324), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n886), .B2(new_n889), .ZN(G1353gat));
  INV_X1    g689(.A(G211gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(KEYINPUT124), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n630), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n869), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT63), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n873), .A2(new_n891), .A3(new_n630), .ZN(new_n898));
  OAI221_X1 g697(.A(new_n893), .B1(KEYINPUT124), .B2(new_n892), .C1(new_n894), .C2(new_n869), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G1354gat));
  NAND3_X1  g699(.A1(new_n871), .A2(new_n271), .A3(new_n872), .ZN(new_n901));
  INV_X1    g700(.A(G218gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n271), .A2(G218gat), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT125), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n879), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n903), .B(KEYINPUT126), .C1(new_n879), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1355gat));
endmodule


