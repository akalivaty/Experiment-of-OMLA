

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  XNOR2_X1 U326 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U327 ( .A(n459), .B(n458), .ZN(n507) );
  XOR2_X1 U328 ( .A(n403), .B(n402), .Z(n525) );
  XOR2_X1 U329 ( .A(G120GAT), .B(G78GAT), .Z(n294) );
  XNOR2_X1 U330 ( .A(n476), .B(n475), .ZN(n532) );
  INV_X1 U331 ( .A(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U332 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U333 ( .A(n404), .B(n294), .ZN(n303) );
  XNOR2_X1 U334 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n475) );
  INV_X1 U335 ( .A(KEYINPUT93), .ZN(n378) );
  XNOR2_X1 U336 ( .A(n304), .B(n303), .ZN(n308) );
  NOR2_X1 U337 ( .A1(n521), .A2(n434), .ZN(n548) );
  XNOR2_X1 U338 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n386) );
  NOR2_X1 U340 ( .A1(n525), .A2(n482), .ZN(n569) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n460) );
  XNOR2_X1 U342 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U343 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U344 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  INV_X1 U346 ( .A(KEYINPUT73), .ZN(n295) );
  NAND2_X1 U347 ( .A1(n295), .A2(G92GAT), .ZN(n298) );
  INV_X1 U348 ( .A(G92GAT), .ZN(n296) );
  NAND2_X1 U349 ( .A1(n296), .A2(KEYINPUT73), .ZN(n297) );
  NAND2_X1 U350 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n336) );
  XNOR2_X1 U353 ( .A(KEYINPUT76), .B(n336), .ZN(n302) );
  AND2_X1 U354 ( .A1(G230GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n304) );
  XOR2_X1 U356 ( .A(G106GAT), .B(G148GAT), .Z(n404) );
  XOR2_X1 U357 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n306) );
  XNOR2_X1 U358 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U360 ( .A(n308), .B(n307), .Z(n314) );
  XOR2_X1 U361 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n310) );
  XNOR2_X1 U362 ( .A(G71GAT), .B(G57GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n449) );
  XOR2_X1 U364 ( .A(G64GAT), .B(KEYINPUT75), .Z(n312) );
  XNOR2_X1 U365 ( .A(G176GAT), .B(G204GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n371) );
  XNOR2_X1 U367 ( .A(n449), .B(n371), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n580) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G197GAT), .Z(n316) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(G36GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U372 ( .A(n317), .B(G15GAT), .Z(n319) );
  XOR2_X1 U373 ( .A(G113GAT), .B(G1GAT), .Z(n352) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(n352), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U376 ( .A(G29GAT), .B(G43GAT), .Z(n321) );
  XNOR2_X1 U377 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n344) );
  XOR2_X1 U379 ( .A(n344), .B(KEYINPUT67), .Z(n323) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U382 ( .A(n325), .B(n324), .Z(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n327) );
  XNOR2_X1 U384 ( .A(G22GAT), .B(KEYINPUT71), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U386 ( .A(G8GAT), .B(KEYINPUT69), .Z(n329) );
  XNOR2_X1 U387 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n574) );
  NOR2_X1 U391 ( .A1(n580), .A2(n574), .ZN(n492) );
  XOR2_X1 U392 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n335) );
  XNOR2_X1 U393 ( .A(KEYINPUT78), .B(KEYINPUT11), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n348) );
  XOR2_X1 U395 ( .A(G50GAT), .B(G162GAT), .Z(n408) );
  XOR2_X1 U396 ( .A(n336), .B(n408), .Z(n338) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U399 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n340) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(G106GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U402 ( .A(n342), .B(n341), .Z(n346) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n343), .B(G218GAT), .ZN(n375) );
  XNOR2_X1 U405 ( .A(n344), .B(n375), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U407 ( .A(n348), .B(n347), .Z(n568) );
  XOR2_X1 U408 ( .A(KEYINPUT36), .B(n568), .Z(n590) );
  XOR2_X1 U409 ( .A(G85GAT), .B(G162GAT), .Z(n350) );
  XNOR2_X1 U410 ( .A(G29GAT), .B(G127GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(n352), .B(n351), .Z(n354) );
  NAND2_X1 U413 ( .A1(G225GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n368) );
  XOR2_X1 U415 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n356) );
  XNOR2_X1 U416 ( .A(KEYINPUT92), .B(G57GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U418 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n358) );
  XNOR2_X1 U419 ( .A(G155GAT), .B(G148GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U421 ( .A(n360), .B(n359), .Z(n366) );
  XOR2_X1 U422 ( .A(G120GAT), .B(KEYINPUT82), .Z(n362) );
  XNOR2_X1 U423 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n395) );
  XOR2_X1 U425 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n364) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n420) );
  XNOR2_X1 U428 ( .A(n395), .B(n420), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n521) );
  XOR2_X1 U431 ( .A(KEYINPUT79), .B(G211GAT), .Z(n370) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(G183GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n448) );
  XNOR2_X1 U434 ( .A(n371), .B(n448), .ZN(n377) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U437 ( .A(G197GAT), .B(KEYINPUT21), .Z(n405) );
  XNOR2_X1 U438 ( .A(n405), .B(G92GAT), .ZN(n379) );
  XOR2_X1 U439 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U442 ( .A(G169GAT), .B(n384), .ZN(n403) );
  INV_X1 U443 ( .A(n403), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n523) );
  INV_X1 U445 ( .A(n523), .ZN(n428) );
  XOR2_X1 U446 ( .A(G176GAT), .B(G99GAT), .Z(n388) );
  XNOR2_X1 U447 ( .A(G43GAT), .B(G190GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U449 ( .A(G183GAT), .B(KEYINPUT83), .Z(n390) );
  XNOR2_X1 U450 ( .A(KEYINPUT87), .B(KEYINPUT85), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U452 ( .A(n392), .B(n391), .Z(n401) );
  XOR2_X1 U453 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n394) );
  XNOR2_X1 U454 ( .A(G113GAT), .B(G71GAT), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n399) );
  XNOR2_X1 U456 ( .A(G15GAT), .B(G127GAT), .ZN(n438) );
  XNOR2_X1 U457 ( .A(n438), .B(n395), .ZN(n397) );
  NAND2_X1 U458 ( .A1(G227GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n402) );
  INV_X1 U462 ( .A(n525), .ZN(n534) );
  NAND2_X1 U463 ( .A1(n428), .A2(n534), .ZN(n423) );
  XOR2_X1 U464 ( .A(G211GAT), .B(G218GAT), .Z(n407) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n409) );
  XOR2_X1 U467 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U468 ( .A(G204GAT), .B(KEYINPUT24), .Z(n411) );
  NAND2_X1 U469 ( .A1(G228GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U471 ( .A(KEYINPUT91), .B(n412), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n416) );
  XNOR2_X1 U474 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U476 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U477 ( .A(G22GAT), .B(G155GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n419), .B(G78GAT), .ZN(n441) );
  XNOR2_X1 U479 ( .A(n420), .B(n441), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n480) );
  NAND2_X1 U481 ( .A1(n423), .A2(n480), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n424), .B(KEYINPUT97), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n425), .B(KEYINPUT25), .ZN(n431) );
  XNOR2_X1 U484 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n427) );
  NOR2_X1 U485 ( .A1(n534), .A2(n480), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n572) );
  XOR2_X1 U487 ( .A(n428), .B(KEYINPUT27), .Z(n434) );
  INV_X1 U488 ( .A(n434), .ZN(n429) );
  NAND2_X1 U489 ( .A1(n572), .A2(n429), .ZN(n430) );
  NAND2_X1 U490 ( .A1(n431), .A2(n430), .ZN(n432) );
  NAND2_X1 U491 ( .A1(n521), .A2(n432), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n433), .B(KEYINPUT98), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n480), .B(KEYINPUT28), .ZN(n528) );
  NAND2_X1 U494 ( .A1(n548), .A2(n528), .ZN(n533) );
  XNOR2_X1 U495 ( .A(KEYINPUT95), .B(n533), .ZN(n435) );
  NAND2_X1 U496 ( .A1(n435), .A2(n525), .ZN(n436) );
  NAND2_X1 U497 ( .A1(n437), .A2(n436), .ZN(n491) );
  XNOR2_X1 U498 ( .A(G1GAT), .B(G64GAT), .ZN(n440) );
  INV_X1 U499 ( .A(n438), .ZN(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n453) );
  XOR2_X1 U501 ( .A(KEYINPUT15), .B(n441), .Z(n443) );
  NAND2_X1 U502 ( .A1(G231GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n445) );
  XNOR2_X1 U505 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U510 ( .A(n453), .B(n452), .Z(n487) );
  NAND2_X1 U511 ( .A1(n491), .A2(n487), .ZN(n454) );
  XOR2_X1 U512 ( .A(KEYINPUT101), .B(n454), .Z(n455) );
  NOR2_X1 U513 ( .A1(n590), .A2(n455), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT37), .B(n456), .Z(n520) );
  NAND2_X1 U515 ( .A1(n492), .A2(n520), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT38), .B(n457), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n507), .A2(n525), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n461) );
  XOR2_X1 U520 ( .A(n487), .B(KEYINPUT110), .Z(n564) );
  INV_X1 U521 ( .A(n574), .ZN(n562) );
  INV_X1 U522 ( .A(KEYINPUT41), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n580), .B(n464), .ZN(n555) );
  NAND2_X1 U524 ( .A1(n562), .A2(n555), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n564), .A2(n467), .ZN(n468) );
  INV_X1 U528 ( .A(n568), .ZN(n488) );
  NAND2_X1 U529 ( .A1(n468), .A2(n488), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT47), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n590), .A2(n487), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT45), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n471), .A2(n574), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n472), .A2(n580), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n532), .A2(n523), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT54), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n521), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n479), .B(KEYINPUT65), .ZN(n573) );
  AND2_X1 U540 ( .A1(n480), .A2(n573), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n569), .A2(n555), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n484) );
  XNOR2_X1 U544 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n483) );
  INV_X1 U545 ( .A(n487), .ZN(n583) );
  NAND2_X1 U546 ( .A1(n583), .A2(n488), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  AND2_X1 U548 ( .A1(n491), .A2(n490), .ZN(n510) );
  NAND2_X1 U549 ( .A1(n492), .A2(n510), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n521), .A2(n499), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(n493), .Z(n494) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n523), .A2(n499), .ZN(n495) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n525), .A2(n499), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n498), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n528), .A2(n499), .ZN(n500) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U561 ( .A1(n521), .A2(n507), .ZN(n505) );
  XOR2_X1 U562 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n502) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(KEYINPUT100), .B(n503), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n523), .A2(n507), .ZN(n506) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U569 ( .A1(n528), .A2(n507), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  AND2_X1 U572 ( .A1(n574), .A2(n555), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n519), .A2(n510), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n521), .A2(n516), .ZN(n511) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n516), .ZN(n513) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n516), .ZN(n515) );
  XOR2_X1 U581 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n527), .ZN(n526) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n533), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT112), .B(n536), .Z(n545) );
  NAND2_X1 U599 ( .A1(n545), .A2(n562), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U602 ( .A1(n555), .A2(n545), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT113), .Z(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n543) );
  NAND2_X1 U607 ( .A1(n545), .A2(n564), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U611 ( .A1(n568), .A2(n545), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n572), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n532), .A2(n549), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n559), .A2(n562), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT116), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT117), .B(n554), .Z(n557) );
  NAND2_X1 U622 ( .A1(n559), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n583), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT119), .Z(n561) );
  NAND2_X1 U627 ( .A1(n559), .A2(n568), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n569), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n569), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT121), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT58), .B(n567), .Z(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n589) );
  NOR2_X1 U639 ( .A1(n574), .A2(n589), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT123), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n589), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT125), .Z(n586) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

