//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT70), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(KEYINPUT70), .B2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(KEYINPUT71), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT68), .B1(new_n476), .B2(G125), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  OAI211_X1 g054(.A(KEYINPUT68), .B(G125), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n475), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n474), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  INV_X1    g063(.A(new_n465), .ZN(new_n489));
  NAND3_X1  g064(.A1(KEYINPUT70), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n463), .B1(new_n489), .B2(new_n490), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G124), .ZN(new_n503));
  OR2_X1    g078(.A1(G100), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n496), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G162));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n464), .B2(new_n465), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n508), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(KEYINPUT4), .B1(new_n476), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n513));
  OR2_X1    g088(.A1(G102), .A2(G2105), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n514), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G164));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n522));
  INV_X1    g097(.A(new_n518), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n522), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n522), .A2(new_n532), .A3(KEYINPUT75), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT76), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT7), .Z(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(G51), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n524), .A2(new_n525), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n543), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n544), .B2(new_n523), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(new_n530), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n518), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n520), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n550), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n530), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n549), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n520), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT78), .ZN(G188));
  NAND2_X1  g142(.A1(new_n530), .A2(G53), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n520), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n527), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  NAND2_X1  g150(.A1(new_n530), .A2(G49), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT79), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n518), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(G87), .A2(new_n527), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n527), .A2(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n530), .A2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n520), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n520), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n530), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n527), .A2(G85), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n595));
  OR3_X1    g170(.A1(new_n549), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n549), .B2(new_n594), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n596), .A2(new_n597), .B1(G54), .B2(new_n530), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n520), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(new_n599), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(new_n560), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n603), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n619));
  INV_X1    g194(.A(G123), .ZN(new_n620));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  OAI221_X1 g196(.A(new_n619), .B1(new_n501), .B2(new_n620), .C1(new_n621), .C2(new_n494), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(G2096), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n476), .A2(new_n468), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(G14), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT84), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n647), .A3(new_n643), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n653), .B(KEYINPUT17), .Z(new_n658));
  OAI211_X1 g233(.A(new_n656), .B(new_n657), .C1(new_n658), .C2(new_n650), .ZN(new_n659));
  INV_X1    g234(.A(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n653), .A2(new_n651), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n650), .A3(new_n660), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  INV_X1    g259(.A(new_n682), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n679), .A2(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n667), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n683), .A2(new_n687), .A3(new_n667), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  NAND2_X1  g267(.A1(new_n476), .A2(G127), .ZN(new_n693));
  INV_X1    g268(.A(G115), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n467), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n463), .B1(new_n695), .B2(KEYINPUT98), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT98), .B2(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT25), .Z(new_n699));
  INV_X1    g274(.A(G139), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n699), .C1(new_n700), .C2(new_n494), .ZN(new_n701));
  MUX2_X1   g276(.A(G33), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT99), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G2072), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G32), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n495), .A2(G141), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n502), .A2(G129), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT26), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n711), .A2(new_n712), .B1(G105), .B2(new_n468), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n707), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n706), .B1(new_n715), .B2(new_n705), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT27), .ZN(new_n717));
  INV_X1    g292(.A(G1996), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n704), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n604), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G4), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT94), .B(G1348), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n722), .A2(G20), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT23), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1956), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n726), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G168), .A2(new_n722), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n722), .B2(G21), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n722), .A2(G19), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT95), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n560), .B2(new_n722), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1341), .Z(new_n741));
  OAI211_X1 g316(.A(new_n737), .B(new_n741), .C1(new_n705), .C2(new_n622), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n705), .B1(new_n743), .B2(G28), .ZN(new_n745));
  AND2_X1   g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n722), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n722), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n748), .B1(new_n750), .B2(G1961), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G1961), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g327(.A1(G27), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G164), .B2(G29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2078), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n742), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n735), .A2(new_n736), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT100), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n705), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n705), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT29), .B(G2090), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n733), .A2(new_n756), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G104), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n764), .A2(new_n463), .A3(KEYINPUT96), .ZN(new_n765));
  AOI21_X1  g340(.A(KEYINPUT96), .B1(new_n764), .B2(new_n463), .ZN(new_n766));
  OAI221_X1 g341(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT97), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n492), .A2(new_n493), .A3(G140), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n499), .A2(G128), .A3(new_n500), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n705), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n705), .B1(KEYINPUT24), .B2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(KEYINPUT24), .B2(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n487), .B2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G2084), .Z(new_n780));
  NOR4_X1   g355(.A1(new_n721), .A2(new_n763), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n495), .A2(G131), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n502), .A2(G119), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n463), .A2(G107), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n705), .A2(G25), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT87), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT35), .B(G1991), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n722), .B1(G290), .B2(KEYINPUT89), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(KEYINPUT89), .B2(G290), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n722), .A2(G24), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT88), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT90), .B(G1986), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n795), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n722), .A2(G23), .ZN(new_n802));
  INV_X1    g377(.A(G288), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n722), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT91), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT92), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G6), .A2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n586), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  INV_X1    g386(.A(G1981), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n805), .A2(new_n807), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n808), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n722), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n722), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1971), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT34), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n801), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT34), .B1(new_n815), .B2(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n824), .A3(new_n822), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n782), .B1(new_n826), .B2(new_n827), .ZN(G311));
  INV_X1    g403(.A(new_n827), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n824), .B1(new_n821), .B2(new_n822), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n781), .B1(new_n829), .B2(new_n830), .ZN(G150));
  NAND2_X1  g406(.A1(new_n604), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT102), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT38), .Z(new_n834));
  AND2_X1   g409(.A1(new_n518), .A2(G67), .ZN(new_n835));
  AND2_X1   g410(.A1(G80), .A2(G543), .ZN(new_n836));
  OAI21_X1  g411(.A(G651), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT101), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n527), .A2(G93), .B1(new_n530), .B2(G55), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(KEYINPUT101), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n840), .A2(new_n560), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n560), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n834), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n840), .A2(new_n841), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT104), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT103), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n849), .A2(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(new_n506), .B(new_n622), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n487), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n476), .A2(new_n511), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n513), .A2(new_n515), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT106), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(G164), .A2(KEYINPUT106), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n771), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n714), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n714), .ZN(new_n873));
  OAI211_X1 g448(.A(KEYINPUT107), .B(new_n701), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n871), .A4(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n880));
  INV_X1    g455(.A(G142), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n494), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(G130), .B2(new_n502), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n626), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(new_n787), .Z(new_n885));
  AND2_X1   g460(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n878), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n859), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n878), .A2(new_n885), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n858), .B(G160), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n878), .A2(new_n885), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(G395));
  INV_X1    g471(.A(new_n615), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n845), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n604), .A2(G299), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n730), .A2(new_n603), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n730), .B2(new_n603), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n899), .A3(new_n901), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n898), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n898), .B2(new_n908), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  XOR2_X1   g487(.A(G166), .B(G290), .Z(new_n913));
  XNOR2_X1  g488(.A(G305), .B(G288), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n913), .B(new_n914), .Z(new_n915));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n910), .B(new_n916), .C1(new_n898), .C2(new_n908), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n912), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n912), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n850), .A2(new_n607), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  OAI21_X1  g500(.A(G171), .B1(new_n843), .B2(new_n844), .ZN(new_n926));
  INV_X1    g501(.A(new_n844), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(G301), .A3(new_n842), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G286), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n928), .A3(G168), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n925), .B1(new_n932), .B2(new_n904), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n931), .B(new_n930), .C1(new_n906), .C2(new_n909), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n913), .B(new_n914), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n915), .A2(new_n934), .A3(new_n933), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n924), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n935), .A2(new_n936), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n939), .A3(new_n893), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(G397));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n866), .A2(new_n867), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n475), .ZN(new_n953));
  OAI21_X1  g528(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT68), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(new_n956), .B2(new_n480), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n484), .B1(new_n957), .B2(new_n463), .ZN(new_n958));
  INV_X1    g533(.A(new_n473), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT71), .B1(new_n466), .B2(new_n469), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n486), .A2(new_n958), .A3(new_n961), .A4(G40), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(G290), .A2(G1986), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT111), .ZN(new_n965));
  AND2_X1   g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(G1996), .A3(new_n714), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n771), .A2(G2067), .ZN(new_n969));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n768), .A2(new_n970), .A3(new_n769), .A4(new_n770), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(KEYINPUT113), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n963), .B2(new_n972), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n968), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n963), .A2(KEYINPUT112), .A3(new_n718), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n979));
  AND4_X1   g554(.A1(G40), .A2(new_n486), .A3(new_n958), .A4(new_n961), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n951), .A3(new_n950), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n981), .B2(G1996), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n714), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT114), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n973), .B(KEYINPUT113), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n978), .A2(new_n982), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n715), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n968), .ZN(new_n989));
  INV_X1    g564(.A(new_n792), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n787), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n787), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n963), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND4_X1   g568(.A1(new_n967), .A2(new_n984), .A3(new_n989), .A4(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT45), .A4(new_n949), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n949), .B1(new_n512), .B2(new_n516), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n951), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n980), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1971), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(KEYINPUT115), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n949), .C1(new_n512), .C2(new_n516), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n980), .A3(KEYINPUT120), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1009), .B2(new_n962), .ZN(new_n1010));
  INV_X1    g585(.A(new_n996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n1008), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1006), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1000), .B1(new_n1013), .B2(G2090), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT117), .B(G8), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n536), .A2(G8), .A3(new_n537), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n536), .A2(G8), .A3(new_n537), .A4(new_n1019), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1016), .B1(new_n962), .B2(new_n1004), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT118), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(new_n1016), .C1(new_n962), .C2(new_n1004), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G1981), .B1(new_n583), .B2(new_n585), .ZN(new_n1030));
  INV_X1    g605(.A(new_n585), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(new_n812), .A3(new_n581), .A4(new_n582), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT119), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1029), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1041), .B(new_n1046), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n962), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1001), .A2(new_n1008), .A3(new_n1003), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1000), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  AND4_X1   g632(.A1(new_n1024), .A2(new_n1039), .A3(new_n1048), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n980), .A2(new_n1059), .A3(new_n995), .A4(new_n997), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT45), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(G2078), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(new_n980), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n485), .A2(G40), .A3(new_n486), .A4(new_n1050), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1054), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1062), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G171), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n485), .A2(G40), .A3(new_n486), .A4(new_n1065), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n736), .B1(new_n1075), .B2(new_n1063), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT121), .B(G2084), .Z(new_n1077));
  NAND3_X1  g652(.A1(new_n1052), .A2(new_n1054), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1015), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G168), .A2(new_n1015), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(KEYINPUT51), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G8), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT51), .B1(new_n1084), .B2(new_n1080), .ZN(new_n1085));
  AOI211_X1 g660(.A(G168), .B(new_n1015), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1086));
  OAI221_X1 g661(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1082), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1085), .A2(new_n1086), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1058), .A2(new_n1074), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1029), .A2(new_n1037), .A3(new_n1034), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1037), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1041), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1029), .A2(new_n1095), .A3(new_n1045), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1094), .A2(new_n1097), .A3(new_n1057), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n803), .A2(new_n1040), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1032), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1029), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1956), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1013), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n730), .B(KEYINPUT57), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT56), .B(G2072), .Z(new_n1105));
  NOR2_X1   g680(.A1(new_n998), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1348), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n980), .A2(new_n970), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n603), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1104), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1012), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1009), .A2(new_n962), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(KEYINPUT120), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1956), .B1(new_n1117), .B2(new_n1010), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1118), .B2(new_n1106), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT61), .B1(new_n1119), .B2(new_n1108), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n980), .A2(new_n718), .A3(new_n995), .A4(new_n997), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n962), .B2(new_n1004), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n560), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1128), .A3(new_n560), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1348), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n962), .A2(new_n1004), .A3(G2067), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1131), .A2(new_n604), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n1133), .B2(new_n1112), .ZN(new_n1134));
  OR4_X1    g709(.A1(KEYINPUT60), .A2(new_n1131), .A3(new_n603), .A4(new_n1132), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1121), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1119), .A2(new_n1108), .A3(KEYINPUT61), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1120), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1068), .A2(new_n1140), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n961), .A2(G40), .A3(new_n1066), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n463), .B1(new_n482), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1142), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(new_n952), .A3(new_n995), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1141), .A2(G301), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT54), .B1(new_n1148), .B2(new_n1073), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1088), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1056), .A2(G8), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n1023), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1094), .A2(new_n1152), .A3(new_n1097), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(G171), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1072), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(G301), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1072), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1150), .A2(new_n1153), .A3(new_n1024), .A4(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1091), .B(new_n1101), .C1(new_n1139), .C2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1058), .A2(G168), .A3(new_n1079), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1079), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1023), .B2(new_n1151), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1164), .A2(new_n1165), .B1(new_n1153), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n994), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n965), .A2(new_n963), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT125), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n965), .A2(new_n1172), .A3(new_n963), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1175), .A2(new_n984), .A3(new_n989), .A4(new_n993), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT124), .B1(new_n986), .B2(KEYINPUT46), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n978), .A2(new_n982), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n715), .A2(new_n969), .A3(new_n971), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n986), .A2(KEYINPUT46), .B1(new_n963), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1184), .A2(KEYINPUT47), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT47), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1176), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n984), .A2(new_n989), .A3(new_n992), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n981), .B1(new_n1189), .B2(new_n971), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n971), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n963), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1184), .B(KEYINPUT47), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1176), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1169), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g773(.A(G401), .ZN(new_n1200));
  NOR2_X1   g774(.A1(G227), .A2(new_n461), .ZN(new_n1201));
  NAND4_X1  g775(.A1(new_n1200), .A2(KEYINPUT127), .A3(new_n691), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n1203));
  INV_X1    g777(.A(new_n690), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1201), .B1(new_n1204), .B2(new_n688), .ZN(new_n1205));
  OAI21_X1  g779(.A(new_n1203), .B1(new_n1205), .B2(G401), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g781(.A(new_n894), .B(new_n1207), .C1(new_n940), .C2(new_n941), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


