//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  NAND2_X1  g0001(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(KEYINPUT65), .ZN(new_n206));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G50), .ZN(new_n210));
  AOI21_X1  g0010(.A(KEYINPUT65), .B1(new_n210), .B2(new_n207), .ZN(new_n211));
  NOR3_X1   g0011(.A1(new_n209), .A2(new_n211), .A3(G77), .ZN(G353));
  OAI21_X1  g0012(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n208), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n215), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  INV_X1    g0029(.A(G250), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n232));
  INV_X1    g0032(.A(G58), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  INV_X1    g0034(.A(G68), .ZN(new_n235));
  INV_X1    g0035(.A(G238), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n232), .B1(new_n233), .B2(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n217), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n220), .B(new_n225), .C1(KEYINPUT1), .C2(new_n238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n238), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n234), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  INV_X1    g0049(.A(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT66), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n201), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(new_n233), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G223), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n272), .A2(G222), .B1(G77), .B2(new_n271), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n259), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n259), .A3(G274), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n259), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(G179), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n287), .A2(new_n214), .A3(G13), .A4(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n223), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(KEYINPUT70), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n214), .A2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT8), .B(G58), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n215), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(G150), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(KEYINPUT68), .B1(new_n306), .B2(new_n304), .C1(new_n302), .C2(new_n303), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n206), .B1(new_n205), .B2(new_n208), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n207), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n215), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n291), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n286), .A2(new_n288), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n201), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n301), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n283), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n284), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n274), .A2(new_n323), .A3(new_n282), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(KEYINPUT9), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n209), .B2(new_n211), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(new_n309), .A3(new_n310), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n291), .B1(new_n201), .B2(new_n316), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT9), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n301), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(G200), .B2(new_n283), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n325), .A2(new_n330), .ZN(new_n334));
  INV_X1    g0134(.A(new_n324), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT73), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n322), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n283), .A2(G200), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT72), .B(KEYINPUT10), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n321), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n263), .A2(new_n264), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(G20), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n235), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n233), .A2(new_n235), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n207), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n305), .A2(G159), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n345), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT7), .B1(new_n271), .B2(new_n215), .ZN(new_n356));
  NOR4_X1   g0156(.A1(new_n269), .A2(new_n270), .A3(new_n346), .A4(G20), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n354), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n355), .A2(new_n360), .A3(new_n291), .ZN(new_n361));
  INV_X1    g0161(.A(new_n302), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n289), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n302), .B1(new_n214), .B2(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n297), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n259), .A2(G232), .A3(new_n280), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n278), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT76), .ZN(new_n369));
  OR2_X1    g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n279), .A2(G1698), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n371), .C1(new_n269), .C2(new_n270), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n259), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G179), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n278), .A2(new_n367), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n369), .A2(new_n376), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n278), .B2(new_n367), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n259), .B1(new_n372), .B2(new_n373), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(G169), .B1(new_n384), .B2(new_n379), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT18), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n366), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n366), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n369), .A2(new_n376), .A3(new_n323), .A4(new_n379), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n278), .A2(new_n367), .A3(new_n378), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n392), .A2(new_n382), .A3(new_n383), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n393), .B2(G200), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(new_n361), .A3(new_n365), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n396));
  XOR2_X1   g0196(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n266), .A2(G238), .A3(new_n267), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n272), .A2(G232), .B1(G107), .B2(new_n271), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n259), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n278), .B1(new_n228), .B2(new_n281), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n377), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n319), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(new_n293), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(G77), .A3(new_n298), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G20), .A2(G77), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT15), .B(G87), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n303), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n362), .B2(new_n305), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n408), .B1(G77), .B2(new_n289), .C1(new_n292), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n404), .B2(G190), .ZN(new_n415));
  OAI21_X1  g0215(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n390), .A2(new_n399), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n407), .A2(G68), .A3(new_n298), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT12), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n289), .B2(G68), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n316), .A2(KEYINPUT12), .A3(new_n235), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT75), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT75), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n419), .A2(new_n425), .A3(new_n421), .A4(new_n422), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n306), .A2(new_n201), .B1(new_n215), .B2(G68), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n303), .A2(new_n227), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n291), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT11), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(G226), .A2(G1698), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n234), .B2(G1698), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n437), .B2(new_n347), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT74), .B1(new_n438), .B2(new_n259), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n279), .A2(new_n260), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n234), .A2(G1698), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(new_n269), .C2(new_n270), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT74), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(new_n375), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n278), .B1(new_n236), .B2(new_n281), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n433), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(KEYINPUT13), .B(new_n447), .C1(new_n439), .C2(new_n445), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n432), .B(G169), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n444), .B1(new_n443), .B2(new_n375), .ZN(new_n452));
  AOI211_X1 g0252(.A(KEYINPUT74), .B(new_n259), .C1(new_n442), .C2(new_n434), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n446), .A2(new_n433), .A3(new_n448), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(G179), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n432), .B1(new_n459), .B2(G169), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n431), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n424), .A2(new_n426), .A3(new_n430), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(G200), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n463), .C1(new_n323), .C2(new_n459), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n418), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n344), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n228), .A2(G1698), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G238), .B2(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n470), .A2(new_n271), .B1(new_n262), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n375), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n230), .B1(new_n276), .B2(G1), .ZN(new_n474));
  INV_X1    g0274(.A(G274), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n214), .A2(new_n475), .A3(G45), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n259), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n259), .A2(new_n474), .A3(new_n476), .A4(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n323), .ZN(new_n483));
  NOR3_X1   g0283(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT81), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(KEYINPUT19), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT19), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(KEYINPUT81), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n435), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n484), .B1(new_n489), .B2(new_n215), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n215), .A2(G33), .A3(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n215), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT82), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(G20), .B1(new_n263), .B2(new_n264), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G68), .B1(new_n491), .B2(new_n492), .ZN(new_n498));
  INV_X1    g0298(.A(new_n484), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n487), .A2(KEYINPUT81), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n485), .A2(KEYINPUT19), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n434), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n502), .B2(G20), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n496), .A2(new_n291), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n482), .A2(G200), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n214), .A2(G33), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n289), .A2(new_n292), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n316), .A2(new_n410), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n506), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n483), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n498), .A2(new_n503), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n292), .B1(new_n515), .B2(KEYINPUT82), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n505), .B1(new_n316), .B2(new_n410), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n517), .A2(KEYINPUT83), .A3(new_n507), .A4(new_n510), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n375), .A2(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n377), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n482), .A2(new_n319), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n523), .A3(new_n377), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n410), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n509), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n506), .A2(new_n511), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n514), .A2(new_n518), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n289), .A2(G116), .A3(new_n292), .A4(new_n508), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n316), .A2(new_n471), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n290), .A2(new_n223), .B1(G20), .B2(new_n471), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n215), .C1(G33), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT20), .B1(new_n532), .B2(new_n535), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT84), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI211_X1 g0339(.A(KEYINPUT84), .B(KEYINPUT20), .C1(new_n532), .C2(new_n535), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n530), .B(new_n531), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n214), .B(G45), .C1(new_n275), .C2(KEYINPUT5), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT5), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(G41), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n223), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n475), .B1(new_n546), .B2(new_n258), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n260), .A2(G257), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G264), .A2(G1698), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n269), .C2(new_n270), .ZN(new_n551));
  INV_X1    g0351(.A(G303), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n263), .A2(new_n552), .A3(new_n264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n375), .A3(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G270), .B(new_n259), .C1(new_n542), .C2(new_n544), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n548), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n556), .A2(G169), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n541), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n541), .A2(new_n557), .A3(KEYINPUT21), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n548), .A2(new_n554), .A3(G179), .A4(new_n555), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n541), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n556), .A2(new_n323), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n566), .B(new_n541), .C1(G200), .C2(new_n556), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G250), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT78), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(new_n260), .C1(new_n269), .C2(new_n270), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n347), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n533), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n375), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G257), .B(new_n259), .C1(new_n542), .C2(new_n544), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n548), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n377), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n305), .A2(G77), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n582), .A2(new_n534), .A3(G107), .ZN(new_n583));
  XNOR2_X1  g0383(.A(G97), .B(G107), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n581), .B1(new_n585), .B2(new_n215), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n250), .B1(new_n348), .B2(new_n349), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n291), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n316), .A2(new_n534), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n289), .A2(G97), .A3(new_n292), .A4(new_n508), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n571), .A2(new_n572), .B1(G33), .B2(G283), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT78), .B1(new_n265), .B2(G250), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT78), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n569), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n594), .B(new_n574), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n578), .B1(new_n598), .B2(new_n375), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n580), .B(new_n593), .C1(G169), .C2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(G264), .B(new_n259), .C1(new_n542), .C2(new_n544), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G250), .B(new_n260), .C1(new_n269), .C2(new_n270), .ZN(new_n603));
  OAI211_X1 g0403(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G294), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n602), .B1(new_n375), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n377), .A3(new_n548), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n375), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n548), .A3(new_n601), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n319), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n262), .A2(new_n471), .A3(G20), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT23), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n215), .B2(G107), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n250), .A2(KEYINPUT23), .A3(G20), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT22), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n497), .B2(G87), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n215), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(KEYINPUT22), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT24), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(KEYINPUT22), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n347), .A2(new_n617), .A3(new_n215), .A4(G87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT24), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n616), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n292), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n509), .A2(G107), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT25), .B1(new_n289), .B2(G107), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n289), .A2(KEYINPUT25), .A3(G107), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n608), .B(new_n611), .C1(new_n628), .C2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n632), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n625), .A2(new_n626), .A3(new_n616), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n625), .B2(new_n616), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n291), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n610), .A2(G190), .ZN(new_n638));
  AOI21_X1  g0438(.A(G200), .B1(new_n607), .B2(new_n548), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n634), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n576), .A2(G190), .A3(new_n579), .ZN(new_n641));
  OAI21_X1  g0441(.A(G107), .B1(new_n356), .B2(new_n357), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n584), .A2(new_n582), .ZN(new_n643));
  INV_X1    g0443(.A(new_n583), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G20), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(new_n646), .A3(new_n581), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n591), .B1(new_n647), .B2(new_n291), .ZN(new_n648));
  INV_X1    g0448(.A(G200), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n641), .B(new_n648), .C1(new_n649), .C2(new_n599), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n600), .A2(new_n633), .A3(new_n640), .A4(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n468), .A2(new_n529), .A3(new_n568), .A4(new_n651), .ZN(G372));
  INV_X1    g0452(.A(new_n321), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n405), .A2(new_n406), .A3(new_n413), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n464), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n461), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n399), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n390), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n329), .B1(new_n328), .B2(new_n301), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n329), .A2(new_n301), .A3(new_n315), .A4(new_n317), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n332), .B(new_n335), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n339), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n331), .A2(new_n332), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT10), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n341), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n653), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n522), .A2(new_n520), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n528), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  INV_X1    g0470(.A(new_n600), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n640), .A2(new_n650), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n558), .A2(new_n559), .B1(new_n541), .B2(new_n563), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n633), .A2(new_n673), .A3(new_n561), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n512), .A2(new_n483), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n670), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n529), .A2(KEYINPUT26), .A3(new_n671), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n669), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n666), .B1(new_n467), .B2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n214), .A2(new_n215), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n541), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n568), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n565), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(KEYINPUT85), .B(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n633), .A2(new_n640), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n686), .B1(new_n628), .B2(new_n632), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n686), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n633), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n689), .A2(new_n686), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n611), .A2(new_n608), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n637), .B2(new_n634), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(new_n695), .B1(new_n703), .B2(new_n698), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n218), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n499), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n710), .A2(KEYINPUT86), .B1(new_n707), .B2(new_n222), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(KEYINPUT86), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n650), .B(new_n640), .C1(new_n565), .C2(new_n703), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n676), .B1(new_n714), .B2(new_n600), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n678), .B1(new_n715), .B2(KEYINPUT26), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n686), .B1(new_n716), .B2(new_n668), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n506), .A2(new_n511), .A3(new_n527), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n522), .A2(new_n520), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(new_n512), .B2(new_n483), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n672), .A3(new_n600), .A4(new_n674), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n512), .A2(new_n513), .ZN(new_n725));
  INV_X1    g0525(.A(new_n483), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n518), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n525), .A2(new_n528), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n600), .A2(KEYINPUT26), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT26), .B1(new_n722), .B2(new_n600), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT88), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n668), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n724), .A2(new_n730), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n718), .B1(new_n734), .B2(new_n698), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n576), .A2(new_n579), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n563), .A2(new_n519), .A3(new_n607), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n519), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n739), .A2(new_n556), .A3(new_n610), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n609), .A2(new_n601), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n482), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n599), .A2(new_n745), .A3(KEYINPUT30), .A4(new_n563), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n747), .B2(new_n686), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n744), .A2(new_n482), .A3(new_n562), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT30), .B1(new_n749), .B2(new_n599), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n610), .A2(new_n377), .A3(new_n482), .A4(new_n556), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n599), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT87), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT87), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n741), .A2(new_n743), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n753), .A2(new_n746), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n686), .A2(KEYINPUT31), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n748), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n651), .A2(new_n529), .A3(new_n568), .A4(new_n698), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n691), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n737), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n713), .B1(new_n761), .B2(G1), .ZN(G364));
  AND2_X1   g0562(.A1(new_n215), .A2(G13), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n214), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n707), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n694), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n692), .B2(new_n690), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n766), .B(KEYINPUT89), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n218), .A2(new_n347), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT90), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(G355), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n771), .B2(G355), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G116), .B2(new_n218), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n256), .A2(G45), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n347), .B(new_n706), .C1(new_n276), .C2(new_n222), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n223), .B1(G20), .B2(new_n319), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n769), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n323), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT91), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n377), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G159), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT32), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n649), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G107), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n215), .A2(new_n323), .A3(new_n649), .A4(G179), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT92), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT92), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n229), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n323), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n215), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n534), .ZN(new_n800));
  NAND3_X1  g0600(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n323), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n201), .A2(new_n803), .B1(new_n805), .B2(new_n235), .ZN(new_n806));
  NAND2_X1  g0606(.A1(G20), .A2(G179), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n807), .A2(new_n323), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n347), .B1(new_n809), .B2(new_n227), .C1(new_n233), .C2(new_n811), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n797), .A2(new_n800), .A3(new_n806), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n790), .A2(new_n792), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  INV_X1    g0615(.A(G326), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n809), .A2(new_n815), .B1(new_n803), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n799), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G294), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT33), .B(G317), .Z(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n271), .B1(new_n805), .B2(new_n821), .C1(new_n822), .C2(new_n811), .ZN(new_n823));
  INV_X1    g0623(.A(new_n796), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(G303), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n791), .A2(G283), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n788), .A2(G329), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n814), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n784), .B1(new_n829), .B2(new_n781), .ZN(new_n830));
  INV_X1    g0630(.A(new_n780), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n690), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n768), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n654), .A2(new_n698), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n415), .A2(new_n416), .B1(new_n413), .B2(new_n686), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n654), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n417), .A2(new_n414), .A3(new_n698), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n717), .A2(new_n838), .B1(new_n679), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n760), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n766), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  INV_X1    g0643(.A(new_n769), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n781), .A2(new_n778), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n227), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n791), .ZN(new_n847));
  INV_X1    g0647(.A(new_n788), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n229), .A2(new_n847), .B1(new_n848), .B2(new_n815), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n800), .B1(G283), .B2(new_n804), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n552), .B2(new_n803), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n796), .A2(new_n250), .ZN(new_n852));
  INV_X1    g0652(.A(G294), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n271), .B1(new_n809), .B2(new_n471), .C1(new_n853), .C2(new_n811), .ZN(new_n854));
  NOR4_X1   g0654(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n824), .A2(G50), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n788), .A2(G132), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n791), .A2(G68), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n271), .B1(new_n818), .B2(G58), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT94), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G143), .A2(new_n810), .B1(new_n808), .B2(G159), .ZN(new_n862));
  INV_X1    g0662(.A(G137), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n862), .B1(new_n803), .B2(new_n863), .C1(new_n304), .C2(new_n805), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT34), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n855), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n781), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n846), .B1(new_n866), .B2(new_n867), .C1(new_n838), .C2(new_n779), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n843), .A2(new_n868), .ZN(G384));
  OR2_X1    g0669(.A1(new_n645), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n645), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(G116), .A3(new_n224), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OR3_X1    g0674(.A1(new_n221), .A2(new_n227), .A3(new_n351), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n210), .A2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n214), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT70), .B1(new_n289), .B2(new_n292), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n294), .B(new_n291), .C1(new_n286), .C2(new_n288), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n364), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n363), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n358), .A2(new_n359), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n292), .B1(new_n884), .B2(new_n345), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(new_n360), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n380), .B1(new_n393), .B2(G169), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT18), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n366), .A2(new_n386), .A3(new_n387), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n684), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n431), .A2(new_n686), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n461), .A2(new_n464), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n431), .B(new_n686), .C1(new_n458), .C2(new_n460), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n839), .B1(new_n716), .B2(new_n668), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n414), .A2(new_n686), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(new_n684), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n366), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT96), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n394), .A2(new_n361), .A3(new_n365), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n887), .B1(new_n361), .B2(new_n365), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n902), .B(new_n395), .C1(new_n886), .C2(new_n887), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n684), .B1(new_n361), .B2(new_n365), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n910), .B2(KEYINPUT96), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n902), .B1(new_n390), .B2(new_n399), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n899), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT97), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT17), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n886), .B2(new_n394), .ZN(new_n918));
  AND4_X1   g0718(.A1(new_n361), .A2(new_n394), .A3(new_n365), .A4(new_n397), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n910), .B1(new_n920), .B2(new_n890), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n912), .A4(new_n908), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n916), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n913), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n924), .A2(KEYINPUT97), .A3(KEYINPUT38), .A4(new_n921), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n891), .B1(new_n898), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT98), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT98), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n891), .C1(new_n898), .C2(new_n926), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n923), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n909), .B(new_n900), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n899), .B1(new_n932), .B2(new_n914), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n922), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n656), .A2(new_n698), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n928), .A2(new_n930), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n666), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n737), .B2(new_n468), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n940), .B(new_n942), .Z(new_n943));
  AND3_X1   g0743(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n748), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n759), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n946), .A2(new_n838), .A3(new_n895), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n923), .A3(new_n925), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n933), .B2(new_n922), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n895), .A3(new_n838), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT99), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n946), .A2(new_n895), .A3(KEYINPUT99), .A4(new_n838), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n467), .B1(new_n759), .B2(new_n945), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n692), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT100), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(new_n957), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n943), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n214), .B2(new_n763), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n943), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n878), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT101), .ZN(G367));
  NAND2_X1  g0767(.A1(new_n701), .A2(new_n695), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n699), .B2(new_n701), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n694), .B(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n761), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n671), .A2(new_n686), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n600), .B(new_n650), .C1(new_n648), .C2(new_n698), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n704), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n704), .A2(new_n974), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  INV_X1    g0779(.A(new_n700), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n977), .B2(new_n979), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n971), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n761), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n707), .B(KEYINPUT41), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n764), .ZN(new_n987));
  INV_X1    g0787(.A(new_n974), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n968), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT42), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n600), .B1(new_n973), .B2(new_n633), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n698), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT102), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n517), .A2(new_n510), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n686), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n723), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n669), .A2(new_n996), .A3(new_n686), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n999), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n993), .A2(new_n994), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT43), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1005), .A2(new_n1007), .B1(new_n700), .B2(new_n988), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n700), .A2(new_n988), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1004), .C1(new_n1010), .C2(new_n1006), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n987), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT106), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n706), .A2(new_n347), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n247), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n783), .B1(new_n706), .B2(new_n526), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n844), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT104), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n347), .B1(new_n809), .B2(new_n210), .C1(new_n304), .C2(new_n811), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n824), .B2(G58), .ZN(new_n1021));
  INV_X1    g0821(.A(G159), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n805), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n799), .A2(new_n235), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G143), .C2(new_n802), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n791), .A2(G77), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n788), .A2(G137), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n271), .B1(new_n811), .B2(new_n552), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n818), .A2(G107), .B1(new_n802), .B2(G311), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n853), .B2(new_n805), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G283), .C2(new_n808), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n791), .A2(G97), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT105), .B(G317), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1032), .B(new_n1033), .C1(new_n848), .C2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n796), .A2(new_n471), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT46), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1028), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT47), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n867), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1019), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n998), .A2(new_n780), .A3(new_n999), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1013), .A2(new_n1014), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n986), .A2(new_n764), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1044), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT106), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(G387));
  NOR2_X1   g0850(.A1(new_n971), .A2(new_n708), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n761), .B2(new_n970), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1034), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1053), .A2(new_n810), .B1(new_n808), .B2(G303), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n803), .B2(new_n822), .C1(new_n815), .C2(new_n805), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n824), .A2(G294), .B1(G283), .B2(new_n818), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n271), .B1(new_n848), .B2(new_n816), .C1(new_n471), .C2(new_n847), .ZN(new_n1064));
  OR3_X1    g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n802), .A2(G159), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT108), .Z(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n824), .B2(G77), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n347), .B1(new_n811), .B2(new_n201), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n799), .A2(new_n410), .B1(new_n805), .B2(new_n302), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G68), .C2(new_n808), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n788), .A2(G150), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1071), .A3(new_n1033), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n867), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n362), .A2(new_n201), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT50), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n709), .B(new_n276), .C1(new_n235), .C2(new_n227), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1015), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT107), .Z(new_n1079));
  INV_X1    g0879(.A(new_n244), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n276), .B2(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(G107), .B2(new_n218), .C1(new_n709), .C2(new_n770), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n844), .B(new_n1074), .C1(new_n1082), .C2(new_n782), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(KEYINPUT109), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n699), .A2(new_n831), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(KEYINPUT109), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1086), .A2(new_n1087), .B1(new_n765), .B2(new_n970), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1052), .A2(new_n1088), .ZN(G393));
  NAND2_X1  g0889(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(new_n981), .Z(new_n1091));
  OAI211_X1 g0891(.A(new_n707), .B(new_n983), .C1(new_n1091), .C2(new_n971), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n988), .A2(new_n780), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n253), .A2(new_n1015), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n783), .B1(G97), .B2(new_n706), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n844), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT111), .Z(new_n1097));
  NOR2_X1   g0897(.A1(new_n799), .A2(new_n471), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n271), .B1(new_n805), .B2(new_n552), .C1(new_n853), .C2(new_n809), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n824), .C2(G283), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n792), .C1(new_n822), .C2(new_n848), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G311), .A2(new_n810), .B1(new_n802), .B2(G317), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT112), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(KEYINPUT112), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G87), .A2(new_n791), .B1(new_n788), .B2(G143), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G159), .A2(new_n810), .B1(new_n802), .B2(G150), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT51), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n824), .A2(G68), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n799), .A2(new_n227), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n347), .B1(new_n809), .B2(new_n302), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n205), .C2(new_n804), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1105), .A2(new_n1106), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1097), .B1(new_n781), .B2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1091), .A2(new_n765), .B1(new_n1093), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1092), .A2(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(G330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n945), .B2(new_n759), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n838), .A3(new_n895), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n835), .B1(new_n679), .B2(new_n839), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n938), .B1(new_n1123), .B2(new_n895), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n936), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n938), .B1(new_n933), .B2(new_n922), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n836), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n414), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n600), .B(new_n668), .C1(new_n512), .C2(new_n483), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n714), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n698), .B(new_n1129), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1133), .A2(KEYINPUT113), .A3(new_n835), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT113), .B1(new_n1133), .B2(new_n835), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1127), .B1(new_n1136), .B2(new_n895), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1122), .B1(new_n1125), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1133), .A2(new_n835), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT113), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1133), .A2(KEYINPUT113), .A3(new_n835), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n895), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1126), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n760), .A2(new_n838), .A3(new_n895), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n936), .C2(new_n1124), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n895), .B1(new_n1120), .B2(new_n838), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n691), .B(new_n837), .C1(new_n758), .C2(new_n759), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1121), .B1(new_n1152), .B2(new_n895), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1150), .A2(new_n1151), .B1(new_n1123), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n344), .A2(new_n466), .A3(new_n1120), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n735), .B1(new_n717), .B2(new_n718), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n666), .B(new_n1155), .C1(new_n1156), .C2(new_n467), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n708), .B1(new_n1148), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1138), .A2(new_n1147), .A3(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1138), .A2(new_n765), .A3(new_n1147), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n845), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n769), .B1(new_n362), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n271), .B1(new_n811), .B2(new_n471), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1166), .B(new_n797), .C1(G97), .C2(new_n808), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n805), .A2(new_n250), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1168), .B(new_n1111), .C1(G283), .C2(new_n802), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n788), .A2(G294), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n858), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n304), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G125), .B2(new_n788), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n271), .B1(new_n791), .B2(new_n205), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT114), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT53), .B1(new_n796), .B2(new_n304), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1178), .A2(new_n808), .B1(new_n810), .B2(G132), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n803), .B2(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n799), .A2(new_n1022), .B1(new_n805), .B2(new_n863), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1174), .A2(KEYINPUT114), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1171), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1165), .B1(new_n1186), .B2(new_n781), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n936), .B2(new_n779), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1163), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT115), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1163), .A2(KEYINPUT115), .A3(new_n1188), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1162), .A2(new_n1191), .A3(new_n1192), .ZN(G378));
  NAND3_X1  g0993(.A1(new_n950), .A2(G330), .A3(new_n956), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n318), .A2(new_n901), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n665), .B2(new_n321), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n653), .B(new_n1196), .C1(new_n664), .C2(new_n341), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n343), .A2(new_n1196), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1195), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n665), .A2(new_n321), .A3(new_n1197), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1200), .A2(KEYINPUT118), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1194), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n1204), .A3(KEYINPUT118), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1207), .A2(G330), .A3(new_n950), .A4(new_n956), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n940), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n927), .A2(KEYINPUT98), .B1(new_n938), .B2(new_n936), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1211), .A2(new_n1206), .A3(new_n930), .A4(new_n1208), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1157), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1210), .A2(new_n1212), .B1(new_n1161), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n707), .B1(new_n1214), .B2(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1161), .A2(new_n1213), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1216), .A2(new_n1217), .A3(KEYINPUT57), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1200), .A2(new_n1204), .A3(new_n778), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n766), .B1(new_n205), .B2(new_n1164), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(G33), .A2(G41), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT116), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n201), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n275), .B2(new_n271), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n847), .A2(new_n233), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n824), .A2(G77), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n803), .A2(new_n471), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1228), .B(new_n1024), .C1(G97), .C2(new_n804), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n526), .A2(new_n808), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G41), .B(new_n347), .C1(G107), .C2(new_n810), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1226), .B(new_n1232), .C1(G283), .C2(new_n788), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1225), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n811), .A2(new_n1180), .B1(new_n809), .B2(new_n863), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G132), .B2(new_n804), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n818), .A2(G150), .B1(new_n802), .B2(G125), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n796), .C2(new_n1177), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1223), .B1(new_n788), .B2(G124), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n1022), .C2(new_n847), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1235), .B1(new_n1240), .B2(new_n1243), .C1(new_n1234), .C2(new_n1233), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1221), .B1(new_n1244), .B2(new_n781), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1216), .A2(new_n765), .B1(new_n1220), .B2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1219), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1159), .A2(new_n985), .A3(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT119), .Z(new_n1251));
  OAI21_X1  g1051(.A(new_n769), .B1(G68), .B2(new_n1164), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n895), .A2(new_n779), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n824), .A2(G97), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n802), .A2(G294), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n818), .A2(new_n526), .B1(new_n804), .B2(G116), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n809), .A2(new_n250), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n347), .B(new_n1257), .C1(G283), .C2(new_n810), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1026), .B1(new_n848), .B2(new_n552), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n824), .A2(G159), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n802), .A2(G132), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n818), .A2(G50), .B1(new_n804), .B2(new_n1178), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n347), .B1(new_n809), .B2(new_n304), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G137), .B2(new_n810), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n233), .A2(new_n847), .B1(new_n848), .B2(new_n1180), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1259), .A2(new_n1260), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1252), .B(new_n1253), .C1(new_n781), .C2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1154), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n764), .B(KEYINPUT120), .Z(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1269), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1251), .A2(new_n1273), .ZN(G381));
  NOR4_X1   g1074(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G390), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1189), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1278), .A2(G375), .ZN(G407));
  NAND2_X1  g1079(.A1(new_n685), .A2(G213), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT121), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1247), .A2(new_n1277), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G407), .A2(G213), .A3(new_n1282), .ZN(G409));
  XNOR2_X1  g1083(.A(G393), .B(new_n833), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1013), .A2(new_n1044), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1286), .A2(G390), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1276), .B2(new_n1287), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1286), .A2(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(G390), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n1284), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1246), .C1(new_n1215), .C2(new_n1218), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1210), .A2(KEYINPUT122), .A3(new_n1212), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT122), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1271), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1216), .A2(new_n1217), .A3(new_n985), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1220), .A2(new_n1245), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1277), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1281), .B1(new_n1294), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT60), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1249), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT123), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1303), .A2(KEYINPUT123), .A3(new_n1249), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1249), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n708), .B1(new_n1308), .B2(KEYINPUT60), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1310), .A2(G384), .A3(new_n1273), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1310), .B2(new_n1273), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1292), .A2(new_n1293), .A3(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(G2897), .A3(new_n1281), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1281), .A2(G2897), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1302), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1315), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT124), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1294), .A2(new_n1301), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1281), .ZN(new_n1326));
  AND4_X1   g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .A4(new_n1313), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1324), .B1(new_n1302), .B2(new_n1313), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1323), .B1(KEYINPUT63), .B2(new_n1329), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1293), .B1(new_n1331), .B2(new_n1302), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1302), .A2(KEYINPUT62), .A3(new_n1313), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1333), .B1(new_n1335), .B2(KEYINPUT126), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1337), .B(new_n1334), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1332), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1292), .B(KEYINPUT127), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1330), .B1(new_n1339), .B2(new_n1340), .ZN(G405));
  INV_X1    g1141(.A(new_n1277), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1294), .B1(new_n1247), .B2(new_n1342), .ZN(new_n1343));
  XOR2_X1   g1143(.A(new_n1343), .B(new_n1313), .Z(new_n1344));
  XNOR2_X1  g1144(.A(new_n1340), .B(new_n1344), .ZN(G402));
endmodule


