

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(G160), .A2(G40), .ZN(n669) );
  NOR2_X2 U550 ( .A1(G164), .A2(G1384), .ZN(n764) );
  NAND2_X1 U551 ( .A1(n699), .A2(n698), .ZN(n701) );
  AND2_X1 U552 ( .A1(n746), .A2(n988), .ZN(n747) );
  NOR2_X1 U553 ( .A1(n678), .A2(n992), .ZN(n684) );
  XNOR2_X1 U554 ( .A(n715), .B(KEYINPUT94), .ZN(n688) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n700) );
  NOR2_X1 U556 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U557 ( .A(KEYINPUT102), .ZN(n761) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n518), .ZN(n882) );
  XNOR2_X1 U559 ( .A(KEYINPUT15), .B(n569), .ZN(n1007) );
  NOR2_X1 U560 ( .A1(G651), .A2(n621), .ZN(n636) );
  INV_X1 U561 ( .A(G2104), .ZN(n518) );
  NAND2_X1 U562 ( .A1(G101), .A2(n882), .ZN(n514) );
  XOR2_X1 U563 ( .A(KEYINPUT23), .B(n514), .Z(n517) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n515), .Z(n881) );
  NAND2_X1 U566 ( .A1(n881), .A2(G137), .ZN(n516) );
  NAND2_X1 U567 ( .A1(n517), .A2(n516), .ZN(n523) );
  AND2_X1 U568 ( .A1(n518), .A2(G2105), .ZN(n886) );
  NAND2_X1 U569 ( .A1(G125), .A2(n886), .ZN(n521) );
  NAND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XOR2_X1 U571 ( .A(KEYINPUT64), .B(n519), .Z(n889) );
  NAND2_X1 U572 ( .A1(G113), .A2(n889), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U574 ( .A1(n523), .A2(n522), .ZN(G160) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n621) );
  NAND2_X1 U576 ( .A1(G52), .A2(n636), .ZN(n526) );
  INV_X1 U577 ( .A(G651), .ZN(n527) );
  NOR2_X1 U578 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n524), .Z(n637) );
  NAND2_X1 U580 ( .A1(G64), .A2(n637), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U583 ( .A1(G90), .A2(n632), .ZN(n529) );
  NOR2_X2 U584 ( .A1(n621), .A2(n527), .ZN(n633) );
  NAND2_X1 U585 ( .A1(G77), .A2(n633), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(n530), .Z(n531) );
  NOR2_X1 U588 ( .A1(n532), .A2(n531), .ZN(G171) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G57), .ZN(G237) );
  NAND2_X1 U591 ( .A1(G138), .A2(n881), .ZN(n534) );
  NAND2_X1 U592 ( .A1(G102), .A2(n882), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G126), .A2(n886), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G114), .A2(n889), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U597 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U598 ( .A1(n632), .A2(G89), .ZN(n539) );
  XNOR2_X1 U599 ( .A(n539), .B(KEYINPUT4), .ZN(n541) );
  NAND2_X1 U600 ( .A1(G76), .A2(n633), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U602 ( .A(KEYINPUT5), .B(n542), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n637), .A2(G63), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT73), .B(n543), .Z(n545) );
  NAND2_X1 U605 ( .A1(n636), .A2(G51), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n546), .Z(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U609 ( .A(KEYINPUT7), .B(n549), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U613 ( .A(G223), .ZN(n830) );
  NAND2_X1 U614 ( .A1(n830), .A2(G567), .ZN(n551) );
  XOR2_X1 U615 ( .A(KEYINPUT11), .B(n551), .Z(G234) );
  NAND2_X1 U616 ( .A1(G56), .A2(n637), .ZN(n552) );
  XOR2_X1 U617 ( .A(KEYINPUT14), .B(n552), .Z(n558) );
  NAND2_X1 U618 ( .A1(n632), .A2(G81), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT12), .ZN(n555) );
  NAND2_X1 U620 ( .A1(G68), .A2(n633), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT13), .B(n556), .Z(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n636), .A2(G43), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n992) );
  INV_X1 U626 ( .A(G860), .ZN(n605) );
  OR2_X1 U627 ( .A1(n992), .A2(n605), .ZN(G153) );
  XNOR2_X1 U628 ( .A(G171), .B(KEYINPUT69), .ZN(G301) );
  NAND2_X1 U629 ( .A1(G66), .A2(n637), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(KEYINPUT70), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G54), .A2(n636), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G92), .A2(n632), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U634 ( .A1(G79), .A2(n633), .ZN(n564) );
  XNOR2_X1 U635 ( .A(KEYINPUT71), .B(n564), .ZN(n565) );
  NOR2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U638 ( .A1(n1007), .A2(G868), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT72), .B(n570), .Z(n572) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(G284) );
  NAND2_X1 U642 ( .A1(G91), .A2(n632), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G78), .A2(n633), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G53), .A2(n636), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G65), .A2(n637), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT67), .B(n577), .Z(n578) );
  NOR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n997) );
  XOR2_X1 U650 ( .A(n997), .B(KEYINPUT68), .Z(G299) );
  NOR2_X1 U651 ( .A1(G299), .A2(G868), .ZN(n581) );
  INV_X1 U652 ( .A(G868), .ZN(n650) );
  NOR2_X1 U653 ( .A1(G286), .A2(n650), .ZN(n580) );
  NOR2_X1 U654 ( .A1(n581), .A2(n580), .ZN(G297) );
  NAND2_X1 U655 ( .A1(n605), .A2(G559), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n582), .A2(n1007), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U658 ( .A1(G868), .A2(n992), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G868), .A2(n1007), .ZN(n584) );
  NOR2_X1 U660 ( .A1(G559), .A2(n584), .ZN(n585) );
  NOR2_X1 U661 ( .A1(n586), .A2(n585), .ZN(G282) );
  NAND2_X1 U662 ( .A1(G123), .A2(n886), .ZN(n587) );
  XNOR2_X1 U663 ( .A(n587), .B(KEYINPUT18), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n882), .A2(G99), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G135), .A2(n881), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G111), .A2(n889), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n971) );
  XNOR2_X1 U670 ( .A(n971), .B(G2096), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n594), .B(KEYINPUT74), .ZN(n596) );
  INV_X1 U672 ( .A(G2100), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(G156) );
  NAND2_X1 U674 ( .A1(G93), .A2(n632), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G80), .A2(n633), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G55), .A2(n636), .ZN(n600) );
  NAND2_X1 U678 ( .A1(G67), .A2(n637), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U680 ( .A(KEYINPUT75), .B(n601), .Z(n602) );
  OR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n651) );
  XNOR2_X1 U682 ( .A(n651), .B(KEYINPUT76), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G559), .A2(n1007), .ZN(n604) );
  XOR2_X1 U684 ( .A(n992), .B(n604), .Z(n648) );
  NAND2_X1 U685 ( .A1(n648), .A2(n605), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n607), .B(n606), .ZN(G145) );
  NAND2_X1 U687 ( .A1(G61), .A2(n637), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G86), .A2(n632), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n633), .A2(G73), .ZN(n610) );
  XOR2_X1 U691 ( .A(KEYINPUT2), .B(n610), .Z(n611) );
  NOR2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U693 ( .A(KEYINPUT79), .B(n613), .Z(n615) );
  NAND2_X1 U694 ( .A1(n636), .A2(G48), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G305) );
  NAND2_X1 U696 ( .A1(G651), .A2(G74), .ZN(n616) );
  XOR2_X1 U697 ( .A(KEYINPUT77), .B(n616), .Z(n618) );
  NAND2_X1 U698 ( .A1(n636), .A2(G49), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U700 ( .A(KEYINPUT78), .B(n619), .ZN(n620) );
  NOR2_X1 U701 ( .A1(n637), .A2(n620), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n621), .A2(G87), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(G288) );
  NAND2_X1 U704 ( .A1(n637), .A2(G60), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G85), .A2(n632), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G72), .A2(n633), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G47), .A2(n636), .ZN(n626) );
  XNOR2_X1 U709 ( .A(KEYINPUT65), .B(n626), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT66), .ZN(G290) );
  NAND2_X1 U713 ( .A1(G88), .A2(n632), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G75), .A2(n633), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G50), .A2(n636), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G62), .A2(n637), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U719 ( .A1(n641), .A2(n640), .ZN(G166) );
  XOR2_X1 U720 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n642) );
  XNOR2_X1 U721 ( .A(G288), .B(n642), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n643), .B(n651), .ZN(n645) );
  XNOR2_X1 U723 ( .A(G290), .B(G166), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U725 ( .A(G299), .B(n646), .Z(n647) );
  XNOR2_X1 U726 ( .A(G305), .B(n647), .ZN(n897) );
  XOR2_X1 U727 ( .A(n897), .B(n648), .Z(n649) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n653) );
  NOR2_X1 U729 ( .A1(G868), .A2(n651), .ZN(n652) );
  NOR2_X1 U730 ( .A1(n653), .A2(n652), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(KEYINPUT20), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(KEYINPUT81), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n656), .A2(G2090), .ZN(n657) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U738 ( .A1(G132), .A2(G82), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n659), .B(KEYINPUT22), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n660), .B(KEYINPUT82), .ZN(n661) );
  NOR2_X1 U741 ( .A1(G218), .A2(n661), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G96), .A2(n662), .ZN(n834) );
  NAND2_X1 U743 ( .A1(n834), .A2(G2106), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G69), .A2(G120), .ZN(n663) );
  NOR2_X1 U745 ( .A1(G237), .A2(n663), .ZN(n664) );
  NAND2_X1 U746 ( .A1(G108), .A2(n664), .ZN(n835) );
  NAND2_X1 U747 ( .A1(n835), .A2(G567), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n666), .A2(n665), .ZN(n836) );
  NAND2_X1 U749 ( .A1(G483), .A2(G661), .ZN(n667) );
  NOR2_X1 U750 ( .A1(n836), .A2(n667), .ZN(n833) );
  NAND2_X1 U751 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U752 ( .A(G166), .ZN(G303) );
  NAND2_X2 U753 ( .A1(n764), .A2(n669), .ZN(n715) );
  INV_X1 U754 ( .A(G1996), .ZN(n940) );
  OR2_X1 U755 ( .A1(n715), .A2(n940), .ZN(n671) );
  XNOR2_X1 U756 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n672) );
  INV_X1 U757 ( .A(n672), .ZN(n670) );
  NAND2_X1 U758 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U759 ( .A1(n715), .A2(n940), .ZN(n673) );
  NAND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n715), .A2(G1341), .ZN(n676) );
  NAND2_X1 U763 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U764 ( .A1(n1007), .A2(n684), .ZN(n679) );
  XNOR2_X1 U765 ( .A(n679), .B(KEYINPUT98), .ZN(n683) );
  INV_X1 U766 ( .A(n688), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n702), .A2(G2067), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G1348), .A2(n715), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n1007), .A2(n684), .ZN(n685) );
  XNOR2_X1 U772 ( .A(n685), .B(KEYINPUT99), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n694) );
  NAND2_X1 U774 ( .A1(n688), .A2(G1956), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT95), .B(n689), .ZN(n692) );
  NAND2_X1 U776 ( .A1(n702), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U777 ( .A(n690), .B(KEYINPUT27), .ZN(n691) );
  NOR2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n695), .A2(n997), .ZN(n693) );
  NAND2_X1 U780 ( .A1(n694), .A2(n693), .ZN(n699) );
  NOR2_X1 U781 ( .A1(n695), .A2(n997), .ZN(n697) );
  XOR2_X1 U782 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n696) );
  XNOR2_X1 U783 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U784 ( .A(n701), .B(n700), .ZN(n706) );
  XNOR2_X1 U785 ( .A(G1961), .B(KEYINPUT93), .ZN(n909) );
  NAND2_X1 U786 ( .A1(n715), .A2(n909), .ZN(n704) );
  XNOR2_X1 U787 ( .A(G2078), .B(KEYINPUT25), .ZN(n939) );
  NAND2_X1 U788 ( .A1(n939), .A2(n702), .ZN(n703) );
  NAND2_X1 U789 ( .A1(n704), .A2(n703), .ZN(n711) );
  NAND2_X1 U790 ( .A1(n711), .A2(G171), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n728) );
  NAND2_X1 U792 ( .A1(G8), .A2(n715), .ZN(n758) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n758), .ZN(n733) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n715), .ZN(n729) );
  NOR2_X1 U795 ( .A1(n733), .A2(n729), .ZN(n707) );
  NAND2_X1 U796 ( .A1(G8), .A2(n707), .ZN(n709) );
  XNOR2_X1 U797 ( .A(KEYINPUT30), .B(KEYINPUT100), .ZN(n708) );
  XNOR2_X1 U798 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U799 ( .A1(G168), .A2(n710), .ZN(n713) );
  NOR2_X1 U800 ( .A1(G171), .A2(n711), .ZN(n712) );
  NOR2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U802 ( .A(KEYINPUT31), .B(n714), .Z(n727) );
  INV_X1 U803 ( .A(G8), .ZN(n720) );
  NOR2_X1 U804 ( .A1(G1971), .A2(n758), .ZN(n717) );
  NOR2_X1 U805 ( .A1(G2090), .A2(n715), .ZN(n716) );
  NOR2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n718), .A2(G303), .ZN(n719) );
  OR2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n722) );
  AND2_X1 U809 ( .A1(n727), .A2(n722), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n728), .A2(n721), .ZN(n725) );
  INV_X1 U811 ( .A(n722), .ZN(n723) );
  OR2_X1 U812 ( .A1(n723), .A2(G286), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U814 ( .A(KEYINPUT32), .B(n726), .Z(n735) );
  NAND2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U816 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U818 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U819 ( .A(n736), .B(KEYINPUT101), .ZN(n751) );
  NOR2_X1 U820 ( .A1(G1976), .A2(G288), .ZN(n742) );
  NOR2_X1 U821 ( .A1(G1971), .A2(G303), .ZN(n737) );
  NOR2_X1 U822 ( .A1(n742), .A2(n737), .ZN(n1001) );
  INV_X1 U823 ( .A(KEYINPUT33), .ZN(n738) );
  AND2_X1 U824 ( .A1(n1001), .A2(n738), .ZN(n739) );
  NAND2_X1 U825 ( .A1(n751), .A2(n739), .ZN(n748) );
  NAND2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n996) );
  INV_X1 U827 ( .A(n758), .ZN(n740) );
  AND2_X1 U828 ( .A1(n996), .A2(n740), .ZN(n741) );
  NOR2_X1 U829 ( .A1(KEYINPUT33), .A2(n741), .ZN(n745) );
  NAND2_X1 U830 ( .A1(n742), .A2(KEYINPUT33), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n758), .A2(n743), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U833 ( .A(G1981), .B(G305), .Z(n988) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n754) );
  NOR2_X1 U835 ( .A1(G2090), .A2(G303), .ZN(n749) );
  NAND2_X1 U836 ( .A1(G8), .A2(n749), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n752), .A2(n758), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n760) );
  NOR2_X1 U840 ( .A1(G1981), .A2(G305), .ZN(n755) );
  XOR2_X1 U841 ( .A(n755), .B(KEYINPUT92), .Z(n756) );
  XNOR2_X1 U842 ( .A(KEYINPUT24), .B(n756), .ZN(n757) );
  NOR2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X2 U844 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U845 ( .A(n762), .B(n761), .ZN(n800) );
  NAND2_X1 U846 ( .A1(G160), .A2(G40), .ZN(n763) );
  NOR2_X1 U847 ( .A1(n764), .A2(n763), .ZN(n815) );
  XNOR2_X1 U848 ( .A(KEYINPUT37), .B(G2067), .ZN(n804) );
  NAND2_X1 U849 ( .A1(G140), .A2(n881), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G104), .A2(n882), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U852 ( .A(KEYINPUT34), .B(n767), .ZN(n774) );
  XNOR2_X1 U853 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n772) );
  NAND2_X1 U854 ( .A1(G116), .A2(n889), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n886), .A2(G128), .ZN(n768) );
  XOR2_X1 U856 ( .A(KEYINPUT83), .B(n768), .Z(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U858 ( .A(n772), .B(n771), .Z(n773) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U860 ( .A(n775), .B(KEYINPUT36), .ZN(n776) );
  XOR2_X1 U861 ( .A(n776), .B(KEYINPUT85), .Z(n864) );
  NOR2_X1 U862 ( .A1(n804), .A2(n864), .ZN(n972) );
  NAND2_X1 U863 ( .A1(n815), .A2(n972), .ZN(n813) );
  NAND2_X1 U864 ( .A1(G141), .A2(n881), .ZN(n777) );
  XNOR2_X1 U865 ( .A(n777), .B(KEYINPUT88), .ZN(n784) );
  NAND2_X1 U866 ( .A1(G129), .A2(n886), .ZN(n779) );
  NAND2_X1 U867 ( .A1(G117), .A2(n889), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n882), .A2(G105), .ZN(n780) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n780), .Z(n781) );
  NOR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U873 ( .A(KEYINPUT89), .B(n785), .ZN(n862) );
  NOR2_X1 U874 ( .A1(n862), .A2(n940), .ZN(n795) );
  NAND2_X1 U875 ( .A1(n889), .A2(G107), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G131), .A2(n881), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G95), .A2(n882), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n886), .A2(G119), .ZN(n788) );
  XOR2_X1 U880 ( .A(KEYINPUT86), .B(n788), .Z(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U883 ( .A(n793), .B(KEYINPUT87), .Z(n863) );
  AND2_X1 U884 ( .A1(n863), .A2(G1991), .ZN(n794) );
  NOR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n964) );
  XOR2_X1 U886 ( .A(n815), .B(KEYINPUT90), .Z(n796) );
  NOR2_X1 U887 ( .A1(n964), .A2(n796), .ZN(n808) );
  INV_X1 U888 ( .A(n808), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n813), .A2(n797), .ZN(n798) );
  XNOR2_X1 U890 ( .A(KEYINPUT91), .B(n798), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U892 ( .A(n801), .B(KEYINPUT103), .ZN(n803) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n1003) );
  NAND2_X1 U894 ( .A1(n1003), .A2(n815), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n818) );
  AND2_X1 U896 ( .A1(n864), .A2(n804), .ZN(n805) );
  XNOR2_X1 U897 ( .A(n805), .B(KEYINPUT105), .ZN(n980) );
  XOR2_X1 U898 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n811) );
  AND2_X1 U899 ( .A1(n940), .A2(n862), .ZN(n961) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n863), .ZN(n970) );
  NOR2_X1 U902 ( .A1(n806), .A2(n970), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n961), .A2(n809), .ZN(n810) );
  XOR2_X1 U905 ( .A(n811), .B(n810), .Z(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n980), .A2(n814), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  XNOR2_X1 U911 ( .A(G2454), .B(G2446), .ZN(n828) );
  XNOR2_X1 U912 ( .A(G2430), .B(G2443), .ZN(n826) );
  XOR2_X1 U913 ( .A(G2435), .B(KEYINPUT106), .Z(n821) );
  XNOR2_X1 U914 ( .A(G2451), .B(G2438), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U916 ( .A(n822), .B(G2427), .Z(n824) );
  XNOR2_X1 U917 ( .A(G1348), .B(G1341), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n824), .B(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n829), .A2(G14), .ZN(n903) );
  XNOR2_X1 U922 ( .A(KEYINPUT107), .B(n903), .ZN(G401) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U925 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U929 ( .A(G132), .ZN(G219) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G82), .ZN(G220) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n836), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2096), .B(G2678), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2072), .B(KEYINPUT43), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n839), .B(KEYINPUT42), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2090), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U942 ( .A(KEYINPUT108), .B(G2100), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1961), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n848), .B(G2474), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1981), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1956), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n886), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n882), .A2(G100), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G136), .A2(n881), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G112), .A2(n889), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U963 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n866) );
  XOR2_X1 U965 ( .A(G164), .B(n864), .Z(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n868) );
  XNOR2_X1 U968 ( .A(G162), .B(KEYINPUT111), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U971 ( .A(G160), .B(n971), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n895) );
  NAND2_X1 U973 ( .A1(G139), .A2(n881), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G103), .A2(n882), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(KEYINPUT110), .B(n875), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G127), .A2(n886), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G115), .A2(n889), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n965) );
  NAND2_X1 U982 ( .A1(G142), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G106), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(KEYINPUT45), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G130), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G118), .A2(n889), .ZN(n890) );
  XNOR2_X1 U989 ( .A(KEYINPUT109), .B(n890), .ZN(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n965), .B(n893), .Z(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n992), .B(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(G171), .B(n1007), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(G286), .B(n900), .Z(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(n902) );
  XNOR2_X1 U999 ( .A(KEYINPUT112), .B(n902), .ZN(G397) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n903), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G96), .ZN(G221) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1009 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n1018) );
  XOR2_X1 U1010 ( .A(G16), .B(KEYINPUT121), .Z(n934) );
  XNOR2_X1 U1011 ( .A(G5), .B(n909), .ZN(n931) );
  XOR2_X1 U1012 ( .A(G1966), .B(G21), .Z(n920) );
  XOR2_X1 U1013 ( .A(G1341), .B(G19), .Z(n913) );
  XNOR2_X1 U1014 ( .A(G1956), .B(G20), .ZN(n911) );
  XNOR2_X1 U1015 ( .A(G1981), .B(G6), .ZN(n910) );
  NOR2_X1 U1016 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1018 ( .A(KEYINPUT122), .B(n914), .ZN(n917) );
  XOR2_X1 U1019 ( .A(KEYINPUT59), .B(G1348), .Z(n915) );
  XNOR2_X1 U1020 ( .A(G4), .B(n915), .ZN(n916) );
  NOR2_X1 U1021 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1022 ( .A(KEYINPUT60), .B(n918), .ZN(n919) );
  NAND2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n921) );
  XNOR2_X1 U1025 ( .A(n921), .B(KEYINPUT58), .ZN(n927) );
  XOR2_X1 U1026 ( .A(G1986), .B(G24), .Z(n925) );
  XNOR2_X1 U1027 ( .A(G1971), .B(G22), .ZN(n923) );
  XNOR2_X1 U1028 ( .A(G23), .B(G1976), .ZN(n922) );
  NOR2_X1 U1029 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1030 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1031 ( .A(n927), .B(n926), .Z(n928) );
  NOR2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(n932), .B(KEYINPUT61), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT125), .B(n935), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n936), .A2(G11), .ZN(n987) );
  XOR2_X1 U1038 ( .A(G2090), .B(G35), .Z(n953) );
  XOR2_X1 U1039 ( .A(G1991), .B(G25), .Z(n937) );
  NAND2_X1 U1040 ( .A1(n937), .A2(G28), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n938), .B(KEYINPUT114), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n939), .B(G27), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(n940), .B(G32), .ZN(n941) );
  NAND2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(KEYINPUT115), .B(n943), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n950), .Z(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT116), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(G34), .B(G2084), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n954), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1057 ( .A(KEYINPUT117), .B(n957), .Z(n958) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n959), .B(KEYINPUT55), .ZN(n985) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n960) );
  NOR2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1062 ( .A(KEYINPUT51), .B(n962), .Z(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n979) );
  XOR2_X1 U1064 ( .A(G2072), .B(n965), .Z(n967) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n968), .ZN(n977) );
  XOR2_X1 U1068 ( .A(G160), .B(G2084), .Z(n969) );
  NOR2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT113), .B(n975), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT52), .B(n982), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(G29), .A2(n983), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n1016) );
  XNOR2_X1 U1080 ( .A(KEYINPUT56), .B(G16), .ZN(n1013) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(KEYINPUT57), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT118), .B(n991), .ZN(n1011) );
  XOR2_X1 U1085 ( .A(G171), .B(G1961), .Z(n994) );
  XNOR2_X1 U1086 ( .A(n992), .B(G1341), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1006) );
  NAND2_X1 U1088 ( .A1(G1971), .A2(G303), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1090 ( .A(n997), .B(G1956), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(KEYINPUT119), .B(n1004), .Z(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(G1348), .B(n1007), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1014), .B(KEYINPUT120), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1018), .B(n1017), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1019), .ZN(G150) );
  INV_X1 U1104 ( .A(G150), .ZN(G311) );
endmodule

