

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U550 ( .A1(n521), .A2(G2104), .ZN(n897) );
  NAND2_X2 U551 ( .A1(n733), .A2(G8), .ZN(n735) );
  INV_X1 U552 ( .A(KEYINPUT64), .ZN(n692) );
  NAND2_X1 U553 ( .A1(n691), .A2(n799), .ZN(n693) );
  NOR2_X1 U554 ( .A1(G1966), .A2(n735), .ZN(n748) );
  XNOR2_X1 U555 ( .A(n743), .B(KEYINPUT32), .ZN(n744) );
  AND2_X1 U556 ( .A1(n742), .A2(n741), .ZN(n745) );
  INV_X1 U557 ( .A(KEYINPUT101), .ZN(n743) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n799) );
  NOR2_X1 U559 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n532), .Z(n652) );
  NOR2_X2 U561 ( .A1(n525), .A2(n524), .ZN(G160) );
  XOR2_X1 U562 ( .A(KEYINPUT29), .B(n714), .Z(n514) );
  AND2_X1 U563 ( .A1(G8), .A2(n747), .ZN(n515) );
  OR2_X1 U564 ( .A1(n701), .A2(n700), .ZN(n704) );
  XNOR2_X1 U565 ( .A(KEYINPUT98), .B(KEYINPUT30), .ZN(n722) );
  XNOR2_X1 U566 ( .A(n723), .B(n722), .ZN(n724) );
  INV_X1 U567 ( .A(KEYINPUT102), .ZN(n760) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n729) );
  INV_X1 U569 ( .A(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U570 ( .A1(n769), .A2(n768), .ZN(n770) );
  INV_X1 U571 ( .A(n820), .ZN(n810) );
  INV_X1 U572 ( .A(KEYINPUT75), .ZN(n595) );
  AND2_X1 U573 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U574 ( .A(n595), .B(KEYINPUT15), .ZN(n596) );
  NOR2_X1 U575 ( .A1(n647), .A2(n537), .ZN(n650) );
  INV_X1 U576 ( .A(KEYINPUT17), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n597), .B(n596), .ZN(n1005) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n647) );
  NAND2_X1 U579 ( .A1(n895), .A2(G137), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n551), .A2(n550), .ZN(G171) );
  NOR2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XNOR2_X2 U582 ( .A(n517), .B(n516), .ZN(n895) );
  INV_X1 U583 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U584 ( .A1(G101), .A2(n897), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n525) );
  NOR2_X2 U587 ( .A1(G2104), .A2(n521), .ZN(n904) );
  NAND2_X1 U588 ( .A1(G125), .A2(n904), .ZN(n523) );
  AND2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U590 ( .A1(G113), .A2(n901), .ZN(n522) );
  NAND2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  AND2_X1 U592 ( .A1(G138), .A2(n895), .ZN(n531) );
  NAND2_X1 U593 ( .A1(G102), .A2(n897), .ZN(n529) );
  NAND2_X1 U594 ( .A1(G126), .A2(n904), .ZN(n527) );
  NAND2_X1 U595 ( .A1(G114), .A2(n901), .ZN(n526) );
  AND2_X1 U596 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(G164) );
  INV_X1 U599 ( .A(G651), .ZN(n537) );
  NOR2_X1 U600 ( .A1(G543), .A2(n537), .ZN(n532) );
  NAND2_X1 U601 ( .A1(G65), .A2(n652), .ZN(n535) );
  NOR2_X1 U602 ( .A1(G651), .A2(n647), .ZN(n533) );
  XNOR2_X2 U603 ( .A(KEYINPUT66), .B(n533), .ZN(n653) );
  NAND2_X1 U604 ( .A1(G53), .A2(n653), .ZN(n534) );
  NAND2_X1 U605 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U606 ( .A(KEYINPUT71), .B(n536), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n650), .A2(G78), .ZN(n538) );
  XOR2_X1 U608 ( .A(KEYINPUT69), .B(n538), .Z(n540) );
  NOR2_X1 U609 ( .A1(G651), .A2(G543), .ZN(n656) );
  NAND2_X1 U610 ( .A1(n656), .A2(G91), .ZN(n539) );
  NAND2_X1 U611 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U612 ( .A(KEYINPUT70), .B(n541), .Z(n542) );
  NAND2_X1 U613 ( .A1(n543), .A2(n542), .ZN(G299) );
  NAND2_X1 U614 ( .A1(G52), .A2(n653), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n652), .A2(G64), .ZN(n544) );
  NAND2_X1 U616 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U617 ( .A1(G90), .A2(n656), .ZN(n547) );
  NAND2_X1 U618 ( .A1(G77), .A2(n650), .ZN(n546) );
  NAND2_X1 U619 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U620 ( .A(KEYINPUT68), .B(n548), .Z(n549) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(n549), .ZN(n550) );
  XOR2_X1 U622 ( .A(G2438), .B(G2454), .Z(n553) );
  XNOR2_X1 U623 ( .A(G2435), .B(G2430), .ZN(n552) );
  XNOR2_X1 U624 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U625 ( .A(n554), .B(G2427), .Z(n556) );
  XNOR2_X1 U626 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U627 ( .A(n556), .B(n555), .ZN(n560) );
  XOR2_X1 U628 ( .A(G2443), .B(G2446), .Z(n558) );
  XNOR2_X1 U629 ( .A(KEYINPUT106), .B(G2451), .ZN(n557) );
  XNOR2_X1 U630 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U631 ( .A(n560), .B(n559), .Z(n561) );
  AND2_X1 U632 ( .A1(G14), .A2(n561), .ZN(G401) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  INV_X1 U635 ( .A(G57), .ZN(G237) );
  NAND2_X1 U636 ( .A1(G89), .A2(n656), .ZN(n562) );
  XNOR2_X1 U637 ( .A(n562), .B(KEYINPUT4), .ZN(n563) );
  XNOR2_X1 U638 ( .A(KEYINPUT76), .B(n563), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n650), .A2(G76), .ZN(n564) );
  XOR2_X1 U640 ( .A(KEYINPUT77), .B(n564), .Z(n565) );
  NAND2_X1 U641 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U642 ( .A(KEYINPUT5), .B(n567), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G63), .A2(n652), .ZN(n569) );
  NAND2_X1 U644 ( .A1(G51), .A2(n653), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n571) );
  XOR2_X1 U646 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n570) );
  XNOR2_X1 U647 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U649 ( .A(KEYINPUT7), .B(n574), .ZN(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U652 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U653 ( .A(G223), .ZN(n830) );
  NAND2_X1 U654 ( .A1(n830), .A2(G567), .ZN(n576) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U656 ( .A1(n656), .A2(G81), .ZN(n577) );
  XNOR2_X1 U657 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U658 ( .A1(G68), .A2(n650), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(n580), .Z(n584) );
  NAND2_X1 U661 ( .A1(G56), .A2(n652), .ZN(n581) );
  XNOR2_X1 U662 ( .A(n581), .B(KEYINPUT73), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n582), .B(KEYINPUT14), .ZN(n583) );
  NOR2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U665 ( .A1(G43), .A2(n653), .ZN(n585) );
  NAND2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n1000) );
  INV_X1 U667 ( .A(n1000), .ZN(n587) );
  NAND2_X1 U668 ( .A1(n587), .A2(G860), .ZN(G153) );
  INV_X1 U669 ( .A(G171), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n650), .A2(G79), .ZN(n589) );
  NAND2_X1 U672 ( .A1(G54), .A2(n653), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U674 ( .A(n590), .B(KEYINPUT74), .ZN(n594) );
  NAND2_X1 U675 ( .A1(G66), .A2(n652), .ZN(n592) );
  NAND2_X1 U676 ( .A1(G92), .A2(n656), .ZN(n591) );
  NAND2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n597) );
  INV_X1 U679 ( .A(G868), .ZN(n671) );
  NAND2_X1 U680 ( .A1(n1005), .A2(n671), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(G284) );
  NOR2_X1 U682 ( .A1(G286), .A2(n671), .ZN(n601) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U684 ( .A1(n601), .A2(n600), .ZN(G297) );
  INV_X1 U685 ( .A(G559), .ZN(n602) );
  NOR2_X1 U686 ( .A1(G860), .A2(n602), .ZN(n603) );
  XNOR2_X1 U687 ( .A(KEYINPUT79), .B(n603), .ZN(n604) );
  INV_X1 U688 ( .A(n1005), .ZN(n839) );
  NAND2_X1 U689 ( .A1(n604), .A2(n839), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(n1005), .A2(n671), .ZN(n606) );
  XOR2_X1 U692 ( .A(KEYINPUT80), .B(n606), .Z(n607) );
  NOR2_X1 U693 ( .A1(G559), .A2(n607), .ZN(n609) );
  NOR2_X1 U694 ( .A1(G868), .A2(n1000), .ZN(n608) );
  NOR2_X1 U695 ( .A1(n609), .A2(n608), .ZN(G282) );
  XOR2_X1 U696 ( .A(G2100), .B(KEYINPUT82), .Z(n619) );
  NAND2_X1 U697 ( .A1(G123), .A2(n904), .ZN(n610) );
  XOR2_X1 U698 ( .A(KEYINPUT81), .B(n610), .Z(n611) );
  XNOR2_X1 U699 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U700 ( .A1(G99), .A2(n897), .ZN(n612) );
  NAND2_X1 U701 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U702 ( .A1(G135), .A2(n895), .ZN(n615) );
  NAND2_X1 U703 ( .A1(G111), .A2(n901), .ZN(n614) );
  NAND2_X1 U704 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U705 ( .A1(n617), .A2(n616), .ZN(n929) );
  XNOR2_X1 U706 ( .A(G2096), .B(n929), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U708 ( .A1(G93), .A2(n656), .ZN(n621) );
  NAND2_X1 U709 ( .A1(G80), .A2(n650), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n652), .A2(G67), .ZN(n622) );
  XNOR2_X1 U712 ( .A(n622), .B(KEYINPUT84), .ZN(n624) );
  NAND2_X1 U713 ( .A1(G55), .A2(n653), .ZN(n623) );
  NAND2_X1 U714 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n672) );
  NAND2_X1 U716 ( .A1(G559), .A2(n839), .ZN(n627) );
  XOR2_X1 U717 ( .A(n1000), .B(n627), .Z(n669) );
  XNOR2_X1 U718 ( .A(KEYINPUT83), .B(n669), .ZN(n628) );
  NOR2_X1 U719 ( .A1(G860), .A2(n628), .ZN(n629) );
  XOR2_X1 U720 ( .A(n672), .B(n629), .Z(G145) );
  NAND2_X1 U721 ( .A1(G85), .A2(n656), .ZN(n631) );
  NAND2_X1 U722 ( .A1(G72), .A2(n650), .ZN(n630) );
  NAND2_X1 U723 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U724 ( .A1(G47), .A2(n653), .ZN(n632) );
  XNOR2_X1 U725 ( .A(KEYINPUT67), .B(n632), .ZN(n633) );
  NOR2_X1 U726 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U727 ( .A1(n652), .A2(G60), .ZN(n635) );
  NAND2_X1 U728 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G61), .A2(n652), .ZN(n638) );
  NAND2_X1 U730 ( .A1(G86), .A2(n656), .ZN(n637) );
  NAND2_X1 U731 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U732 ( .A1(n650), .A2(G73), .ZN(n639) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U734 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U735 ( .A1(G48), .A2(n653), .ZN(n642) );
  NAND2_X1 U736 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U737 ( .A1(G651), .A2(G74), .ZN(n645) );
  NAND2_X1 U738 ( .A1(G49), .A2(n653), .ZN(n644) );
  NAND2_X1 U739 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U740 ( .A1(n652), .A2(n646), .ZN(n649) );
  NAND2_X1 U741 ( .A1(n647), .A2(G87), .ZN(n648) );
  NAND2_X1 U742 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U743 ( .A1(G75), .A2(n650), .ZN(n651) );
  XNOR2_X1 U744 ( .A(n651), .B(KEYINPUT86), .ZN(n661) );
  NAND2_X1 U745 ( .A1(G62), .A2(n652), .ZN(n655) );
  NAND2_X1 U746 ( .A1(G50), .A2(n653), .ZN(n654) );
  NAND2_X1 U747 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U748 ( .A1(G88), .A2(n656), .ZN(n657) );
  XNOR2_X1 U749 ( .A(KEYINPUT85), .B(n657), .ZN(n658) );
  NOR2_X1 U750 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U751 ( .A1(n661), .A2(n660), .ZN(G303) );
  INV_X1 U752 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U753 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U754 ( .A(G288), .B(KEYINPUT88), .ZN(n662) );
  XNOR2_X1 U755 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U756 ( .A(G305), .B(n664), .ZN(n666) );
  INV_X1 U757 ( .A(G299), .ZN(n997) );
  XNOR2_X1 U758 ( .A(n997), .B(G166), .ZN(n665) );
  XNOR2_X1 U759 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U760 ( .A(n672), .B(n667), .ZN(n668) );
  XNOR2_X1 U761 ( .A(G290), .B(n668), .ZN(n840) );
  XOR2_X1 U762 ( .A(n669), .B(n840), .Z(n670) );
  NOR2_X1 U763 ( .A1(n671), .A2(n670), .ZN(n674) );
  NOR2_X1 U764 ( .A1(G868), .A2(n672), .ZN(n673) );
  NOR2_X1 U765 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U766 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U767 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U768 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U769 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U770 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XOR2_X1 U771 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  XNOR2_X1 U772 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U773 ( .A1(G120), .A2(G69), .ZN(n679) );
  NOR2_X1 U774 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U775 ( .A1(G108), .A2(n680), .ZN(n837) );
  NAND2_X1 U776 ( .A1(G567), .A2(n837), .ZN(n687) );
  NOR2_X1 U777 ( .A1(G219), .A2(G220), .ZN(n682) );
  XNOR2_X1 U778 ( .A(KEYINPUT89), .B(KEYINPUT22), .ZN(n681) );
  XNOR2_X1 U779 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U780 ( .A1(n683), .A2(G218), .ZN(n684) );
  XNOR2_X1 U781 ( .A(KEYINPUT90), .B(n684), .ZN(n685) );
  NAND2_X1 U782 ( .A1(n685), .A2(G96), .ZN(n836) );
  NAND2_X1 U783 ( .A1(G2106), .A2(n836), .ZN(n686) );
  NAND2_X1 U784 ( .A1(n687), .A2(n686), .ZN(n917) );
  NAND2_X1 U785 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U786 ( .A1(n917), .A2(n688), .ZN(n835) );
  NAND2_X1 U787 ( .A1(n835), .A2(G36), .ZN(G176) );
  NOR2_X1 U788 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U789 ( .A1(G8), .A2(n689), .ZN(n690) );
  XNOR2_X1 U790 ( .A(n690), .B(KEYINPUT104), .ZN(n751) );
  NAND2_X1 U791 ( .A1(G160), .A2(G40), .ZN(n798) );
  INV_X1 U792 ( .A(n798), .ZN(n691) );
  XNOR2_X2 U793 ( .A(n693), .B(n692), .ZN(n716) );
  NAND2_X1 U794 ( .A1(n716), .A2(G1996), .ZN(n694) );
  XNOR2_X1 U795 ( .A(n694), .B(KEYINPUT26), .ZN(n696) );
  INV_X1 U796 ( .A(n716), .ZN(n733) );
  NAND2_X1 U797 ( .A1(n733), .A2(G1341), .ZN(n695) );
  NAND2_X1 U798 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U799 ( .A1(n1000), .A2(n697), .ZN(n701) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n716), .ZN(n699) );
  NAND2_X1 U801 ( .A1(n733), .A2(G1348), .ZN(n698) );
  NAND2_X1 U802 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U803 ( .A1(n1005), .A2(n702), .ZN(n700) );
  NAND2_X1 U804 ( .A1(n1005), .A2(n702), .ZN(n703) );
  NAND2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n716), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U807 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  AND2_X1 U808 ( .A1(n733), .A2(G1956), .ZN(n706) );
  NOR2_X1 U809 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U810 ( .A1(n997), .A2(n710), .ZN(n708) );
  NAND2_X1 U811 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U812 ( .A1(n997), .A2(n710), .ZN(n711) );
  XOR2_X1 U813 ( .A(n711), .B(KEYINPUT28), .Z(n712) );
  NAND2_X1 U814 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U815 ( .A1(G1961), .A2(n716), .ZN(n715) );
  XNOR2_X1 U816 ( .A(n715), .B(KEYINPUT97), .ZN(n718) );
  XNOR2_X1 U817 ( .A(KEYINPUT25), .B(G2078), .ZN(n976) );
  NAND2_X1 U818 ( .A1(n976), .A2(n716), .ZN(n717) );
  NAND2_X1 U819 ( .A1(n718), .A2(n717), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n725), .A2(G171), .ZN(n719) );
  NAND2_X1 U821 ( .A1(n514), .A2(n719), .ZN(n732) );
  NOR2_X1 U822 ( .A1(n733), .A2(G2084), .ZN(n747) );
  INV_X1 U823 ( .A(n747), .ZN(n720) );
  NAND2_X1 U824 ( .A1(G8), .A2(n720), .ZN(n721) );
  OR2_X1 U825 ( .A1(n748), .A2(n721), .ZN(n723) );
  NOR2_X1 U826 ( .A1(G168), .A2(n724), .ZN(n728) );
  NOR2_X1 U827 ( .A1(G171), .A2(n725), .ZN(n726) );
  XOR2_X1 U828 ( .A(KEYINPUT99), .B(n726), .Z(n727) );
  NOR2_X1 U829 ( .A1(n728), .A2(n727), .ZN(n730) );
  XNOR2_X1 U830 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U831 ( .A1(n732), .A2(n731), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n746), .A2(G286), .ZN(n742) );
  INV_X1 U833 ( .A(G8), .ZN(n740) );
  NOR2_X1 U834 ( .A1(n733), .A2(G2090), .ZN(n734) );
  XNOR2_X1 U835 ( .A(n734), .B(KEYINPUT100), .ZN(n737) );
  NOR2_X1 U836 ( .A1(n735), .A2(G1971), .ZN(n736) );
  NOR2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U838 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U839 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U840 ( .A(n745), .B(n744), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n748), .A2(n515), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n746), .A2(n749), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n755), .A2(n753), .ZN(n750) );
  NAND2_X1 U844 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n752), .A2(n735), .ZN(n778) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  AND2_X1 U847 ( .A1(n753), .A2(n1003), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n759) );
  INV_X1 U849 ( .A(n1003), .ZN(n757) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U852 ( .A1(n766), .A2(n756), .ZN(n1012) );
  OR2_X1 U853 ( .A1(n757), .A2(n1012), .ZN(n758) );
  NAND2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n761) );
  XNOR2_X1 U855 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U856 ( .A1(n735), .A2(n762), .ZN(n763) );
  XNOR2_X1 U857 ( .A(n763), .B(KEYINPUT65), .ZN(n765) );
  AND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n767), .A2(n735), .ZN(n768) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n994) );
  NAND2_X1 U862 ( .A1(n770), .A2(n994), .ZN(n771) );
  XNOR2_X1 U863 ( .A(n771), .B(KEYINPUT103), .ZN(n776) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U865 ( .A(n772), .B(KEYINPUT96), .Z(n773) );
  XNOR2_X1 U866 ( .A(KEYINPUT24), .B(n773), .ZN(n774) );
  NOR2_X1 U867 ( .A1(n735), .A2(n774), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n814) );
  NAND2_X1 U869 ( .A1(G119), .A2(n904), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G107), .A2(n901), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G95), .A2(n897), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G131), .A2(n895), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT91), .B(n783), .Z(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U877 ( .A(KEYINPUT92), .B(n786), .Z(n892) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n892), .ZN(n797) );
  XOR2_X1 U879 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n788) );
  NAND2_X1 U880 ( .A1(G105), .A2(n897), .ZN(n787) );
  XNOR2_X1 U881 ( .A(n788), .B(n787), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G129), .A2(n904), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G117), .A2(n901), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT93), .B(n791), .Z(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n895), .A2(G141), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n875) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n875), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n930) );
  NOR2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n824) );
  NAND2_X1 U892 ( .A1(n930), .A2(n824), .ZN(n800) );
  XNOR2_X1 U893 ( .A(n800), .B(KEYINPUT95), .ZN(n817) );
  NAND2_X1 U894 ( .A1(G104), .A2(n897), .ZN(n802) );
  NAND2_X1 U895 ( .A1(G140), .A2(n895), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n803), .ZN(n808) );
  NAND2_X1 U898 ( .A1(G128), .A2(n904), .ZN(n805) );
  NAND2_X1 U899 ( .A1(G116), .A2(n901), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n806), .Z(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n809), .ZN(n894) );
  XNOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NOR2_X1 U905 ( .A1(n894), .A2(n822), .ZN(n935) );
  NAND2_X1 U906 ( .A1(n935), .A2(n824), .ZN(n820) );
  NOR2_X1 U907 ( .A1(n817), .A2(n810), .ZN(n812) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n1011) );
  NAND2_X1 U909 ( .A1(n1011), .A2(n824), .ZN(n811) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n827) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n875), .ZN(n919) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n892), .ZN(n931) );
  NOR2_X1 U914 ( .A1(n815), .A2(n931), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n919), .A2(n818), .ZN(n819) );
  XNOR2_X1 U917 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n894), .A2(n822), .ZN(n938) );
  NAND2_X1 U920 ( .A1(n823), .A2(n938), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n829) );
  XOR2_X1 U923 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n828) );
  XNOR2_X1 U924 ( .A(n829), .B(n828), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n830), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n832) );
  INV_X1 U927 ( .A(G661), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U932 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  XOR2_X1 U935 ( .A(KEYINPUT109), .B(n838), .Z(G325) );
  XOR2_X1 U936 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U939 ( .A(n839), .B(G286), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n843) );
  XOR2_X1 U941 ( .A(n1000), .B(G171), .Z(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  NOR2_X1 U943 ( .A1(G37), .A2(n844), .ZN(G397) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2084), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n847), .B(G2096), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U950 ( .A(G2100), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U951 ( .A(KEYINPUT111), .B(G2678), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U953 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U954 ( .A(KEYINPUT112), .B(G1991), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1956), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n856), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1971), .B(G1976), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U960 ( .A(G1986), .B(G1981), .Z(n860) );
  XNOR2_X1 U961 ( .A(G1966), .B(G1961), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U964 ( .A(KEYINPUT113), .B(G2474), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U966 ( .A1(n904), .A2(G124), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G136), .A2(n895), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT114), .B(n868), .Z(n870) );
  NAND2_X1 U971 ( .A1(n901), .A2(G112), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G100), .A2(n897), .ZN(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT115), .B(n871), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U976 ( .A(G164), .B(G162), .Z(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U978 ( .A(n876), .B(KEYINPUT48), .Z(n878) );
  XNOR2_X1 U979 ( .A(KEYINPUT120), .B(KEYINPUT46), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(n879), .B(n929), .Z(n890) );
  NAND2_X1 U982 ( .A1(n901), .A2(G115), .ZN(n880) );
  XOR2_X1 U983 ( .A(KEYINPUT119), .B(n880), .Z(n882) );
  NAND2_X1 U984 ( .A1(n904), .A2(G127), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n883), .B(KEYINPUT47), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G139), .A2(n895), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n897), .A2(G103), .ZN(n886) );
  XOR2_X1 U990 ( .A(KEYINPUT118), .B(n886), .Z(n887) );
  NOR2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n922) );
  XNOR2_X1 U992 ( .A(G160), .B(n922), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n909) );
  NAND2_X1 U996 ( .A1(n895), .A2(G142), .ZN(n896) );
  XOR2_X1 U997 ( .A(KEYINPUT117), .B(n896), .Z(n899) );
  NAND2_X1 U998 ( .A1(n897), .A2(G106), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(KEYINPUT45), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n901), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(n904), .A2(G130), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT116), .B(n905), .Z(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n910), .ZN(G395) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n912), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n917), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(KEYINPUT121), .B(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(n914), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n917), .ZN(G319) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(KEYINPUT55), .ZN(n986) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1021 ( .A(KEYINPUT123), .B(n920), .Z(n921) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n921), .Z(n927) );
  XOR2_X1 U1023 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n925), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n940) );
  XOR2_X1 U1028 ( .A(G2084), .B(G160), .Z(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n936), .B(KEYINPUT122), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n986), .A2(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n993) );
  XNOR2_X1 U1039 ( .A(KEYINPUT126), .B(KEYINPUT60), .ZN(n953) );
  XNOR2_X1 U1040 ( .A(KEYINPUT59), .B(G1348), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(G4), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G1956), .B(G20), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1341), .B(G19), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G6), .B(G1981), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(KEYINPUT125), .B(n947), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n953), .B(n952), .ZN(n965) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n957) );
  XNOR2_X1 U1051 ( .A(G1971), .B(G22), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(G23), .B(G1976), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n959), .B(n958), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G21), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G1961), .B(G5), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1062 ( .A(KEYINPUT61), .B(n966), .Z(n967) );
  NOR2_X1 U1063 ( .A1(G16), .A2(n967), .ZN(n991) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G1996), .B(G32), .Z(n970) );
  NAND2_X1 U1069 ( .A1(n970), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(G25), .B(G1991), .ZN(n971) );
  XNOR2_X1 U1071 ( .A(KEYINPUT124), .B(n971), .ZN(n972) );
  NOR2_X1 U1072 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1074 ( .A(G27), .B(n976), .Z(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1078 ( .A(G2084), .B(G34), .Z(n982) );
  XNOR2_X1 U1079 ( .A(KEYINPUT54), .B(n982), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(n986), .B(n985), .ZN(n988) );
  INV_X1 U1082 ( .A(G29), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(G11), .A2(n989), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1019) );
  XOR2_X1 U1087 ( .A(G16), .B(KEYINPUT56), .Z(n1017) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G168), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(n996), .B(KEYINPUT57), .ZN(n1009) );
  XNOR2_X1 U1091 ( .A(n997), .B(G1956), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(G1971), .A2(G303), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(G1341), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G1348), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G301), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(n1020), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

