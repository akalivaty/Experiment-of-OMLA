//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n438, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(new_n438), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT68), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND3_X1   g038(.A1(KEYINPUT70), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(KEYINPUT70), .B2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n468), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT71), .ZN(G160));
  NOR2_X1   g053(.A1(new_n466), .A2(new_n469), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n470), .A2(new_n486), .A3(G138), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n469), .C1(new_n464), .C2(new_n465), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n488), .A2(new_n469), .B1(KEYINPUT4), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n474), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(new_n469), .B2(G114), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(KEYINPUT72), .A3(new_n495), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n491), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n490), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n509), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT73), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n506), .A2(new_n510), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  INV_X1    g096(.A(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT74), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n508), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n511), .A2(new_n531), .B1(new_n513), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n530), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  AOI22_X1  g110(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n508), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT75), .B(G81), .Z(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n511), .A2(new_n538), .B1(new_n513), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  XOR2_X1   g119(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n545));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(G188));
  NOR2_X1   g123(.A1(new_n506), .A2(KEYINPUT79), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT79), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n553));
  AND2_X1   g128(.A1(G78), .A2(G543), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n555), .A2(G651), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n522), .A2(KEYINPUT77), .A3(KEYINPUT9), .A4(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n511), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n522), .A2(G53), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT77), .B(KEYINPUT9), .Z(new_n562));
  AOI22_X1  g137(.A1(new_n560), .A2(G91), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n558), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n560), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n503), .A2(new_n505), .ZN(new_n567));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n508), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n522), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G288));
  NOR2_X1   g146(.A1(new_n520), .A2(KEYINPUT78), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n511), .A2(new_n559), .ZN(new_n573));
  OAI21_X1  g148(.A(G86), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n567), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n578), .A2(new_n579), .B1(G48), .B2(new_n522), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n574), .A2(new_n580), .A3(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n508), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n511), .A2(new_n586), .B1(new_n513), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n560), .A2(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n549), .A2(new_n551), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n593), .B1(G651), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n522), .A2(G54), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n541), .ZN(new_n611));
  MUX2_X1   g186(.A(new_n610), .B(new_n611), .S(KEYINPUT82), .Z(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n479), .A2(G123), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT83), .Z(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(KEYINPUT84), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(KEYINPUT84), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n617), .B(new_n618), .C1(G111), .C2(new_n469), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n467), .A2(G135), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n470), .A2(new_n475), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n622), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2435), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2438), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n633), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(G14), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT88), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n649), .B(KEYINPUT17), .Z(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n647), .A3(new_n645), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n648), .A2(new_n649), .A3(new_n645), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n626), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n665), .A2(KEYINPUT20), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n661), .A3(new_n664), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n670), .C1(KEYINPUT20), .C2(new_n665), .ZN(new_n671));
  XOR2_X1   g246(.A(G1991), .B(G1996), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(G26), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n479), .A2(G128), .ZN(new_n680));
  INV_X1    g255(.A(new_n467), .ZN(new_n681));
  INV_X1    g256(.A(G140), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n684));
  INV_X1    g259(.A(G104), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n469), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT93), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n679), .B1(new_n689), .B2(G29), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n679), .B(new_n690), .S(KEYINPUT28), .Z(new_n691));
  INV_X1    g266(.A(G2067), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G4), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n600), .B2(new_n694), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1348), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n479), .A2(G129), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT98), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT26), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G29), .B2(G32), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT27), .B(G1996), .Z(new_n709));
  AOI21_X1  g284(.A(new_n697), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT30), .B(G28), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G21), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G168), .B2(G16), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G1966), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n694), .A2(G5), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G171), .B2(new_n694), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n712), .B(new_n715), .C1(G1961), .C2(new_n717), .ZN(new_n718));
  OAI22_X1  g293(.A1(new_n717), .A2(G1961), .B1(new_n621), .B2(new_n678), .ZN(new_n719));
  INV_X1    g294(.A(new_n709), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n707), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n714), .A2(G1966), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n718), .A2(new_n721), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(G29), .A2(G33), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n475), .A2(G103), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n467), .A2(G139), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(new_n469), .C2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT95), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(new_n678), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT99), .B1(new_n737), .B2(G29), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n737), .A2(KEYINPUT99), .A3(G29), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n738), .B(new_n739), .C1(G162), .C2(new_n678), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT100), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(G2090), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n694), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n541), .B2(new_n694), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1341), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n724), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n678), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n678), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n710), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G160), .A2(G29), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n756), .A3(new_n678), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2084), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT97), .Z(new_n761));
  OAI21_X1  g336(.A(KEYINPUT23), .B1(new_n604), .B2(new_n694), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n694), .A2(G20), .ZN(new_n763));
  MUX2_X1   g338(.A(KEYINPUT23), .B(new_n762), .S(new_n763), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1956), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n691), .A2(new_n692), .B1(new_n734), .B2(new_n735), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n742), .B2(G2090), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G2084), .B2(new_n759), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n752), .A2(new_n761), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n678), .A2(G25), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n771));
  INV_X1    g346(.A(G131), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n681), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n467), .A2(KEYINPUT89), .A3(G131), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(G119), .B2(new_n479), .ZN(new_n775));
  OR2_X1    g350(.A1(G95), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n770), .B1(new_n778), .B2(new_n678), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT35), .B(G1991), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n694), .A2(G24), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n589), .B2(new_n694), .ZN(new_n783));
  INV_X1    g358(.A(G1986), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n694), .A2(G6), .ZN(new_n786));
  INV_X1    g361(.A(G305), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n694), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n694), .A2(G23), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G288), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT90), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n694), .A2(G22), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n694), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G1971), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n792), .A2(new_n794), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(G1971), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n795), .A2(new_n798), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n790), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n781), .B(new_n785), .C1(new_n802), .C2(KEYINPUT34), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT91), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT92), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n808), .A2(KEYINPUT92), .A3(new_n806), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(KEYINPUT92), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n804), .A2(new_n810), .A3(new_n805), .A4(new_n807), .ZN(new_n811));
  AND4_X1   g386(.A1(new_n693), .A2(new_n769), .A3(new_n809), .A4(new_n811), .ZN(G311));
  NAND4_X1  g387(.A1(new_n769), .A2(new_n809), .A3(new_n693), .A4(new_n811), .ZN(G150));
  AOI22_X1  g388(.A1(new_n520), .A2(G93), .B1(new_n522), .B2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n508), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT37), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n600), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n816), .B(new_n541), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT39), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT101), .Z(G145));
  XNOR2_X1  g401(.A(G160), .B(new_n621), .ZN(new_n827));
  INV_X1    g402(.A(G142), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n681), .A2(KEYINPUT103), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(G106), .A2(G2105), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT103), .B1(new_n681), .B2(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n479), .A2(G130), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n829), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n827), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n704), .B(new_n484), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n500), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT72), .B1(new_n498), .B2(new_n495), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n493), .A2(G2105), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n496), .A2(new_n842), .A3(new_n492), .A4(G2104), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n844), .A2(KEYINPUT102), .A3(new_n491), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n490), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n733), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n688), .ZN(new_n848));
  INV_X1    g423(.A(new_n624), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n778), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n778), .B1(new_n850), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n838), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n848), .B(new_n849), .ZN(new_n857));
  INV_X1    g432(.A(new_n778), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n852), .A3(new_n837), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n855), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g437(.A1(new_n816), .A2(G868), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n864));
  XNOR2_X1  g439(.A(G288), .B(G303), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(G290), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(G290), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n787), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n787), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(KEYINPUT104), .A3(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n869), .A2(KEYINPUT42), .A3(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n600), .A2(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n598), .A2(new_n599), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n604), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n609), .B(new_n821), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n884), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n876), .A2(KEYINPUT105), .A3(new_n877), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n880), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n878), .B(new_n879), .C1(new_n890), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n863), .B1(new_n897), .B2(G868), .ZN(G295));
  AOI21_X1  g473(.A(new_n863), .B1(new_n897), .B2(G868), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n821), .B(G301), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G286), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n886), .A2(new_n887), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n891), .A2(new_n903), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n874), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n874), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n901), .B1(new_n909), .B2(new_n856), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n875), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n905), .A2(new_n874), .A3(new_n906), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n856), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n900), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n901), .A3(new_n856), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT44), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(G397));
  NAND2_X1  g495(.A1(new_n840), .A2(new_n845), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(G2105), .B2(new_n487), .ZN(new_n923));
  AOI21_X1  g498(.A(G1384), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT106), .B(G40), .Z(new_n925));
  NAND2_X1  g500(.A1(new_n477), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n924), .A2(new_n926), .A3(KEYINPUT45), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n778), .A2(new_n780), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n778), .A2(new_n780), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n928), .A2(G1996), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT107), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n688), .B(new_n692), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n704), .B2(G1996), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n933), .A2(new_n704), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n589), .B(new_n784), .ZN(new_n937));
  AOI211_X1 g512(.A(new_n931), .B(new_n936), .C1(new_n927), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n846), .A2(new_n940), .A3(G1384), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n844), .A2(KEYINPUT102), .A3(new_n491), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT102), .B1(new_n844), .B2(new_n491), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n923), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n939), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G2084), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n945), .B1(new_n490), .B2(new_n500), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n926), .B1(KEYINPUT50), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT114), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n940), .B1(new_n846), .B2(G1384), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(KEYINPUT108), .A3(new_n945), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n477), .A2(new_n925), .ZN(new_n957));
  INV_X1    g532(.A(new_n949), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1966), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n947), .A2(new_n963), .A3(new_n948), .A4(new_n950), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G8), .ZN(new_n966));
  NAND2_X1  g541(.A1(G286), .A2(G8), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(KEYINPUT119), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(KEYINPUT51), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(G8), .A3(G286), .ZN(new_n972));
  OAI211_X1 g547(.A(G8), .B(new_n969), .C1(new_n965), .C2(G286), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT50), .B1(new_n953), .B2(new_n955), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n957), .B1(new_n958), .B2(new_n939), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(G2090), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n926), .B1(new_n924), .B2(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n949), .A2(new_n954), .ZN(new_n983));
  AOI21_X1  g558(.A(G1971), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(G8), .B(new_n978), .C1(new_n981), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  INV_X1    g561(.A(new_n984), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n953), .A2(KEYINPUT50), .A3(new_n955), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n958), .A2(new_n939), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n957), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n986), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n985), .B1(new_n992), .B2(new_n978), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT110), .B(G1981), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n574), .A2(new_n580), .A3(new_n582), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n522), .A2(G48), .ZN(new_n997));
  INV_X1    g572(.A(G86), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n581), .C1(new_n998), .C2(new_n511), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G1981), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT111), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT49), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n926), .B1(new_n953), .B2(new_n955), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n986), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n957), .B1(new_n941), .B2(new_n946), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT109), .B1(new_n1006), .B2(G8), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G288), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1009), .A2(G1976), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1004), .B1(new_n1003), .B2(new_n986), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(KEYINPUT109), .A3(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1009), .B2(G1976), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1010), .B(new_n1016), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n994), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n1019), .B2(new_n1010), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1016), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1020), .A2(new_n1022), .A3(KEYINPUT113), .A4(new_n1008), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n993), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n982), .A2(new_n750), .A3(new_n983), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1961), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n979), .B2(new_n980), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n956), .A2(new_n957), .A3(new_n959), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1032), .A2(G171), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n971), .A2(new_n1034), .A3(new_n972), .A4(new_n973), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n975), .A2(new_n1024), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(KEYINPUT122), .A3(new_n1024), .A4(new_n975), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n981), .B2(new_n984), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n977), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1020), .A2(new_n1043), .A3(new_n1022), .A4(new_n1008), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n965), .A2(G8), .A3(G168), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT63), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OR3_X1    g621(.A1(new_n1015), .A2(new_n1017), .A3(new_n985), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT112), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(KEYINPUT112), .ZN(new_n1050));
  AOI211_X1 g625(.A(G1976), .B(G288), .C1(new_n1048), .C2(new_n1002), .ZN(new_n1051));
  INV_X1    g626(.A(new_n996), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1049), .B(new_n1050), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1047), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n965), .A2(new_n1055), .A3(G8), .A4(G168), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n993), .B(new_n1056), .C1(new_n1018), .C2(new_n1023), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G299), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n557), .A2(KEYINPUT57), .A3(new_n558), .A4(new_n563), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n988), .A2(new_n957), .A3(new_n990), .ZN(new_n1063));
  INV_X1    g638(.A(G1956), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n982), .A2(KEYINPUT115), .A3(new_n1066), .A4(new_n983), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n944), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n957), .A3(new_n1066), .A4(new_n983), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1062), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1003), .A2(new_n692), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n979), .A2(new_n980), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(G1348), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT116), .B(new_n1075), .C1(new_n1076), .C2(G1348), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1065), .A2(new_n1072), .A3(new_n1062), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n600), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1074), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1996), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1068), .A2(new_n957), .A3(new_n1085), .A4(new_n983), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT58), .B(G1341), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1003), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT117), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n1086), .C1(new_n1003), .C2(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n541), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1089), .A2(new_n1094), .A3(new_n541), .A4(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1065), .A2(new_n1072), .A3(new_n1062), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT118), .B(new_n1097), .C1(new_n1098), .C2(new_n1073), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1098), .B2(new_n1073), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1082), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT118), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n882), .B1(new_n1081), .B2(KEYINPUT60), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1106), .B(new_n600), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1105), .A2(new_n1107), .B1(KEYINPUT60), .B2(new_n1081), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1084), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(G40), .B1(new_n924), .B2(KEYINPUT45), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1068), .A2(new_n477), .A3(new_n1030), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1027), .B(new_n1029), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1027), .A2(new_n1029), .A3(G301), .A4(new_n1031), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(KEYINPUT54), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1112), .A2(G171), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(new_n1033), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1117), .A2(new_n974), .A3(new_n1024), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1058), .B1(new_n1109), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n938), .B1(new_n1041), .B2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n934), .A2(new_n704), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT46), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1124), .A2(new_n927), .B1(KEYINPUT125), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n933), .B1(new_n1127), .B2(KEYINPUT46), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT107), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n932), .B(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(KEYINPUT125), .A3(new_n1125), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1133), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(new_n1126), .C1(new_n1128), .C2(new_n1131), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n929), .B(KEYINPUT123), .Z(new_n1139));
  OAI221_X1 g714(.A(new_n1138), .B1(G2067), .B2(new_n689), .C1(new_n936), .C2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n935), .A2(new_n928), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1141), .B(new_n1139), .C1(new_n1130), .C2(new_n705), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n689), .A2(G2067), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT124), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1144), .A3(new_n927), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n927), .A2(new_n784), .A3(new_n589), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT48), .Z(new_n1147));
  OR3_X1    g722(.A1(new_n936), .A2(new_n931), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1137), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1137), .A2(new_n1145), .A3(new_n1148), .A4(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1123), .A2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g729(.A1(new_n917), .A2(new_n918), .ZN(new_n1156));
  NOR2_X1   g730(.A1(G229), .A2(new_n462), .ZN(new_n1157));
  AND2_X1   g731(.A1(new_n861), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g732(.A1(G401), .A2(G227), .ZN(new_n1159));
  AND3_X1   g733(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(G308));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(G225));
endmodule


