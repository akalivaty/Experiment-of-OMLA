

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U550 ( .A1(n782), .A2(n776), .ZN(n775) );
  NOR2_X2 U551 ( .A1(n570), .A2(n569), .ZN(G164) );
  NOR2_X1 U552 ( .A1(n800), .A2(n806), .ZN(n516) );
  XOR2_X1 U553 ( .A(n765), .B(n764), .Z(n517) );
  OR2_X1 U554 ( .A1(n783), .A2(n775), .ZN(n778) );
  OR2_X1 U555 ( .A1(n726), .A2(n757), .ZN(n806) );
  XNOR2_X1 U556 ( .A(n691), .B(KEYINPUT65), .ZN(n725) );
  INV_X1 U557 ( .A(n725), .ZN(n693) );
  NOR2_X1 U558 ( .A1(G651), .A2(n641), .ZN(n658) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U560 ( .A1(G85), .A2(n652), .ZN(n519) );
  XOR2_X1 U561 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  INV_X1 U562 ( .A(G651), .ZN(n520) );
  NOR2_X1 U563 ( .A1(n641), .A2(n520), .ZN(n648) );
  NAND2_X1 U564 ( .A1(G72), .A2(n648), .ZN(n518) );
  NAND2_X1 U565 ( .A1(n519), .A2(n518), .ZN(n525) );
  NOR2_X1 U566 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U567 ( .A(KEYINPUT1), .B(n521), .Z(n651) );
  NAND2_X1 U568 ( .A1(G60), .A2(n651), .ZN(n523) );
  NAND2_X1 U569 ( .A1(G47), .A2(n658), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  OR2_X1 U571 ( .A1(n525), .A2(n524), .ZN(G290) );
  XOR2_X1 U572 ( .A(G2438), .B(G2454), .Z(n527) );
  XNOR2_X1 U573 ( .A(G2435), .B(G2430), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U575 ( .A(n528), .B(KEYINPUT108), .Z(n530) );
  XNOR2_X1 U576 ( .A(G1341), .B(G1348), .ZN(n529) );
  XNOR2_X1 U577 ( .A(n530), .B(n529), .ZN(n534) );
  XOR2_X1 U578 ( .A(G2446), .B(G2451), .Z(n532) );
  XNOR2_X1 U579 ( .A(G2443), .B(G2427), .ZN(n531) );
  XNOR2_X1 U580 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U581 ( .A(n534), .B(n533), .Z(n535) );
  AND2_X1 U582 ( .A1(G14), .A2(n535), .ZN(G401) );
  INV_X1 U583 ( .A(G2105), .ZN(n536) );
  AND2_X1 U584 ( .A1(n536), .A2(G2104), .ZN(n884) );
  NAND2_X1 U585 ( .A1(G101), .A2(n884), .ZN(n537) );
  XNOR2_X1 U586 ( .A(n537), .B(KEYINPUT23), .ZN(n538) );
  XNOR2_X1 U587 ( .A(n538), .B(KEYINPUT67), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  XOR2_X2 U589 ( .A(KEYINPUT17), .B(n539), .Z(n885) );
  NAND2_X1 U590 ( .A1(G137), .A2(n885), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n546) );
  NOR2_X1 U592 ( .A1(G2104), .A2(n536), .ZN(n888) );
  NAND2_X1 U593 ( .A1(G125), .A2(n888), .ZN(n544) );
  NAND2_X1 U594 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  XOR2_X2 U595 ( .A(KEYINPUT68), .B(n542), .Z(n890) );
  NAND2_X1 U596 ( .A1(G113), .A2(n890), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U598 ( .A(KEYINPUT66), .B(n547), .ZN(n692) );
  BUF_X1 U599 ( .A(n692), .Z(G160) );
  NAND2_X1 U600 ( .A1(G64), .A2(n651), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G52), .A2(n658), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U603 ( .A1(G90), .A2(n652), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G77), .A2(n648), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U606 ( .A(KEYINPUT9), .B(n552), .ZN(n553) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n553), .ZN(n554) );
  NOR2_X1 U608 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U609 ( .A1(G135), .A2(n885), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G111), .A2(n890), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U612 ( .A1(n888), .A2(G123), .ZN(n558) );
  XOR2_X1 U613 ( .A(KEYINPUT18), .B(n558), .Z(n559) );
  NOR2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U615 ( .A1(n884), .A2(G99), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n918) );
  XNOR2_X1 U617 ( .A(G2096), .B(n918), .ZN(n563) );
  OR2_X1 U618 ( .A1(G2100), .A2(n563), .ZN(G156) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  NAND2_X1 U623 ( .A1(n890), .A2(G114), .ZN(n564) );
  XNOR2_X1 U624 ( .A(n564), .B(KEYINPUT92), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n885), .A2(G138), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G126), .A2(n888), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G102), .A2(n884), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n652), .A2(G89), .ZN(n571) );
  XNOR2_X1 U631 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G76), .A2(n648), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U634 ( .A(n574), .B(KEYINPUT5), .ZN(n579) );
  NAND2_X1 U635 ( .A1(G63), .A2(n651), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G51), .A2(n658), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U638 ( .A(KEYINPUT6), .B(n577), .Z(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U640 ( .A(n580), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G94), .A2(G452), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT70), .B(n581), .Z(G173) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U645 ( .A(n582), .B(KEYINPUT10), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT74), .B(n583), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n833) );
  NAND2_X1 U648 ( .A1(n833), .A2(G567), .ZN(n584) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U650 ( .A1(G56), .A2(n651), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n585), .Z(n591) );
  NAND2_X1 U652 ( .A1(n652), .A2(G81), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G68), .A2(n648), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n589), .Z(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n658), .A2(G43), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n992) );
  XNOR2_X1 U660 ( .A(G860), .B(KEYINPUT75), .ZN(n615) );
  OR2_X1 U661 ( .A1(n992), .A2(n615), .ZN(G153) );
  INV_X1 U662 ( .A(G171), .ZN(G301) );
  NAND2_X1 U663 ( .A1(G66), .A2(n651), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G92), .A2(n652), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G79), .A2(n648), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G54), .A2(n658), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n600), .Z(n601) );
  XNOR2_X1 U671 ( .A(KEYINPUT76), .B(n601), .ZN(n989) );
  INV_X1 U672 ( .A(n989), .ZN(n905) );
  NOR2_X1 U673 ( .A1(n905), .A2(G868), .ZN(n603) );
  INV_X1 U674 ( .A(G868), .ZN(n618) );
  NOR2_X1 U675 ( .A1(n618), .A2(G301), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U677 ( .A1(G91), .A2(n652), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G78), .A2(n648), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT71), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G53), .A2(n658), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n651), .A2(G65), .ZN(n609) );
  XOR2_X1 U684 ( .A(KEYINPUT72), .B(n609), .Z(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U686 ( .A(KEYINPUT73), .B(n612), .ZN(G299) );
  NAND2_X1 U687 ( .A1(G286), .A2(G868), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G299), .A2(n618), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n615), .A2(G559), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n616), .A2(n989), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G559), .A2(n618), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n619), .A2(n989), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n620), .B(KEYINPUT77), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n992), .A2(G868), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G67), .A2(n651), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G55), .A2(n658), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G93), .A2(n652), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G80), .A2(n648), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n665) );
  NAND2_X1 U705 ( .A1(n989), .A2(G559), .ZN(n629) );
  XOR2_X1 U706 ( .A(n992), .B(n629), .Z(n670) );
  XOR2_X1 U707 ( .A(n670), .B(KEYINPUT78), .Z(n630) );
  NOR2_X1 U708 ( .A1(G860), .A2(n630), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT79), .B(n631), .Z(n632) );
  XNOR2_X1 U710 ( .A(n665), .B(n632), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G88), .A2(n652), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT84), .B(n633), .Z(n638) );
  NAND2_X1 U713 ( .A1(G62), .A2(n651), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G50), .A2(n658), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT83), .B(n636), .Z(n637) );
  NOR2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n648), .A2(G75), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(G303) );
  INV_X1 U720 ( .A(G303), .ZN(G166) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U722 ( .A1(G49), .A2(n658), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G87), .A2(n641), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U725 ( .A1(n651), .A2(n644), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n647), .B(KEYINPUT80), .ZN(G288) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n650) );
  NAND2_X1 U729 ( .A1(G73), .A2(n648), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n650), .B(n649), .ZN(n657) );
  NAND2_X1 U731 ( .A1(G61), .A2(n651), .ZN(n654) );
  NAND2_X1 U732 ( .A1(G86), .A2(n652), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U734 ( .A(KEYINPUT81), .B(n655), .Z(n656) );
  NOR2_X1 U735 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n658), .A2(G48), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(G305) );
  NOR2_X1 U738 ( .A1(G868), .A2(n665), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT88), .B(n661), .Z(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n663) );
  XNOR2_X1 U741 ( .A(G166), .B(KEYINPUT85), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(n667) );
  XNOR2_X1 U744 ( .A(G290), .B(G288), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n668), .B(G299), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(G305), .ZN(n904) );
  XNOR2_X1 U748 ( .A(n904), .B(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(G868), .ZN(n672) );
  XOR2_X1 U750 ( .A(KEYINPUT87), .B(n672), .Z(n673) );
  NAND2_X1 U751 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n676), .ZN(n678) );
  XOR2_X1 U755 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n677) );
  XNOR2_X1 U756 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U757 ( .A1(G2072), .A2(n679), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G235), .A2(G236), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT90), .B(n680), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n681), .A2(G57), .ZN(n682) );
  XNOR2_X1 U762 ( .A(KEYINPUT91), .B(n682), .ZN(n683) );
  NAND2_X1 U763 ( .A1(n683), .A2(G108), .ZN(n839) );
  NAND2_X1 U764 ( .A1(G567), .A2(n839), .ZN(n688) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U767 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G96), .A2(n686), .ZN(n840) );
  NAND2_X1 U769 ( .A1(G2106), .A2(n840), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n688), .A2(n687), .ZN(n910) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U772 ( .A1(n910), .A2(n689), .ZN(n838) );
  NAND2_X1 U773 ( .A1(n838), .A2(G36), .ZN(G176) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n691) );
  NAND2_X1 U775 ( .A1(G40), .A2(n692), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n693), .A2(n724), .ZN(n828) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n826) );
  NAND2_X1 U778 ( .A1(G104), .A2(n884), .ZN(n695) );
  NAND2_X1 U779 ( .A1(G140), .A2(n885), .ZN(n694) );
  NAND2_X1 U780 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U781 ( .A(KEYINPUT34), .B(n696), .ZN(n702) );
  NAND2_X1 U782 ( .A1(G128), .A2(n888), .ZN(n698) );
  NAND2_X1 U783 ( .A1(G116), .A2(n890), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U785 ( .A(KEYINPUT93), .B(n699), .ZN(n700) );
  XNOR2_X1 U786 ( .A(KEYINPUT35), .B(n700), .ZN(n701) );
  NOR2_X1 U787 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U788 ( .A(KEYINPUT36), .B(n703), .ZN(n868) );
  NOR2_X1 U789 ( .A1(n826), .A2(n868), .ZN(n928) );
  NAND2_X1 U790 ( .A1(n828), .A2(n928), .ZN(n823) );
  NAND2_X1 U791 ( .A1(G131), .A2(n885), .ZN(n705) );
  NAND2_X1 U792 ( .A1(G107), .A2(n890), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U794 ( .A1(G119), .A2(n888), .ZN(n707) );
  NAND2_X1 U795 ( .A1(G95), .A2(n884), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U798 ( .A(KEYINPUT94), .B(n710), .Z(n867) );
  AND2_X1 U799 ( .A1(G1991), .A2(n867), .ZN(n721) );
  NAND2_X1 U800 ( .A1(G129), .A2(n888), .ZN(n712) );
  NAND2_X1 U801 ( .A1(G117), .A2(n890), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n884), .A2(G105), .ZN(n713) );
  XOR2_X1 U804 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U806 ( .A(KEYINPUT95), .B(n716), .Z(n718) );
  NAND2_X1 U807 ( .A1(n885), .A2(G141), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U809 ( .A(KEYINPUT96), .B(n719), .Z(n901) );
  INV_X1 U810 ( .A(G1996), .ZN(n817) );
  NOR2_X1 U811 ( .A1(n901), .A2(n817), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n926) );
  INV_X1 U813 ( .A(n828), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n926), .A2(n722), .ZN(n820) );
  INV_X1 U815 ( .A(n820), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n823), .A2(n723), .ZN(n809) );
  INV_X1 U817 ( .A(G8), .ZN(n726) );
  NOR2_X2 U818 ( .A1(n725), .A2(n724), .ZN(n757) );
  NOR2_X1 U819 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(KEYINPUT24), .ZN(n728) );
  XNOR2_X1 U821 ( .A(KEYINPUT97), .B(n728), .ZN(n729) );
  OR2_X1 U822 ( .A1(n806), .A2(n729), .ZN(n796) );
  INV_X1 U823 ( .A(G299), .ZN(n1003) );
  INV_X1 U824 ( .A(KEYINPUT98), .ZN(n730) );
  XNOR2_X1 U825 ( .A(n757), .B(n730), .ZN(n756) );
  INV_X1 U826 ( .A(n756), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n742), .A2(G2072), .ZN(n732) );
  XNOR2_X1 U828 ( .A(KEYINPUT100), .B(KEYINPUT27), .ZN(n731) );
  XNOR2_X1 U829 ( .A(n732), .B(n731), .ZN(n734) );
  AND2_X1 U830 ( .A1(n756), .A2(G1956), .ZN(n733) );
  NOR2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n736) );
  NOR2_X1 U832 ( .A1(n1003), .A2(n736), .ZN(n735) );
  XOR2_X1 U833 ( .A(n735), .B(KEYINPUT28), .Z(n753) );
  NAND2_X1 U834 ( .A1(n1003), .A2(n736), .ZN(n751) );
  INV_X1 U835 ( .A(n757), .ZN(n770) );
  NOR2_X1 U836 ( .A1(n770), .A2(n817), .ZN(n737) );
  XOR2_X1 U837 ( .A(n737), .B(KEYINPUT26), .Z(n739) );
  NAND2_X1 U838 ( .A1(n770), .A2(G1341), .ZN(n738) );
  NAND2_X1 U839 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U840 ( .A1(n992), .A2(n740), .ZN(n741) );
  OR2_X1 U841 ( .A1(n989), .A2(n741), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n741), .A2(n989), .ZN(n747) );
  NAND2_X1 U843 ( .A1(G2067), .A2(n742), .ZN(n744) );
  NAND2_X1 U844 ( .A1(G1348), .A2(n770), .ZN(n743) );
  NAND2_X1 U845 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U846 ( .A(KEYINPUT101), .B(n745), .Z(n746) );
  NAND2_X1 U847 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U848 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U849 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U850 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U851 ( .A(KEYINPUT102), .B(KEYINPUT29), .ZN(n754) );
  XNOR2_X1 U852 ( .A(n755), .B(n754), .ZN(n762) );
  XOR2_X1 U853 ( .A(G2078), .B(KEYINPUT25), .Z(n943) );
  NOR2_X1 U854 ( .A1(n943), .A2(n756), .ZN(n759) );
  NOR2_X1 U855 ( .A1(n757), .A2(G1961), .ZN(n758) );
  NOR2_X1 U856 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U857 ( .A(KEYINPUT99), .B(n760), .ZN(n766) );
  AND2_X1 U858 ( .A1(n766), .A2(G171), .ZN(n761) );
  NOR2_X1 U859 ( .A1(n762), .A2(n761), .ZN(n783) );
  XNOR2_X1 U860 ( .A(KEYINPUT30), .B(KEYINPUT103), .ZN(n765) );
  NOR2_X1 U861 ( .A1(G1966), .A2(n806), .ZN(n785) );
  NOR2_X1 U862 ( .A1(G2084), .A2(n770), .ZN(n781) );
  NOR2_X1 U863 ( .A1(n785), .A2(n781), .ZN(n763) );
  NAND2_X1 U864 ( .A1(n763), .A2(G8), .ZN(n764) );
  NOR2_X1 U865 ( .A1(G168), .A2(n517), .ZN(n768) );
  NOR2_X1 U866 ( .A1(G171), .A2(n766), .ZN(n767) );
  NOR2_X1 U867 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U868 ( .A(n769), .B(KEYINPUT31), .ZN(n782) );
  NOR2_X1 U869 ( .A1(G1971), .A2(n806), .ZN(n772) );
  NOR2_X1 U870 ( .A1(G2090), .A2(n770), .ZN(n771) );
  NOR2_X1 U871 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U872 ( .A1(G303), .A2(n773), .ZN(n774) );
  NOR2_X1 U873 ( .A1(n726), .A2(n774), .ZN(n776) );
  OR2_X1 U874 ( .A1(n776), .A2(G286), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n780) );
  XNOR2_X1 U876 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n779) );
  XNOR2_X1 U877 ( .A(n780), .B(n779), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n781), .A2(G8), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G8), .A2(G166), .ZN(n790) );
  NOR2_X1 U884 ( .A1(G2090), .A2(n790), .ZN(n791) );
  XNOR2_X1 U885 ( .A(n791), .B(KEYINPUT105), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n799), .A2(n792), .ZN(n793) );
  XNOR2_X1 U887 ( .A(n793), .B(KEYINPUT106), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n794), .A2(n806), .ZN(n795) );
  AND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X2 U890 ( .A1(n809), .A2(n797), .ZN(n814) );
  NOR2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n804) );
  NOR2_X1 U892 ( .A1(G1971), .A2(G303), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n804), .A2(n798), .ZN(n999) );
  NAND2_X1 U894 ( .A1(n799), .A2(n999), .ZN(n801) );
  NAND2_X1 U895 ( .A1(G1976), .A2(G288), .ZN(n998) );
  INV_X1 U896 ( .A(n998), .ZN(n800) );
  AND2_X1 U897 ( .A1(n801), .A2(n516), .ZN(n802) );
  XNOR2_X1 U898 ( .A(n802), .B(KEYINPUT64), .ZN(n803) );
  NOR2_X1 U899 ( .A1(KEYINPUT33), .A2(n803), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n804), .A2(KEYINPUT33), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n812) );
  XOR2_X1 U903 ( .A(G1981), .B(G305), .Z(n986) );
  INV_X1 U904 ( .A(n809), .ZN(n810) );
  AND2_X1 U905 ( .A1(n986), .A2(n810), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n1006) );
  NAND2_X1 U909 ( .A1(n1006), .A2(n828), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n831) );
  AND2_X1 U911 ( .A1(n817), .A2(n901), .ZN(n921) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n867), .ZN(n917) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n917), .A2(n818), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n921), .A2(n821), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U919 ( .A(KEYINPUT107), .B(n825), .Z(n827) );
  NAND2_X1 U920 ( .A1(n826), .A2(n868), .ZN(n936) );
  NAND2_X1 U921 ( .A1(n827), .A2(n936), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U927 ( .A(G661), .ZN(n834) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n836), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U933 ( .A(G108), .ZN(G238) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G57), .ZN(G237) );
  NOR2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n842) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2072), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1976), .B(G1966), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1971), .B(G1961), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(G1981), .B(G1956), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2474), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U956 ( .A(G1986), .B(KEYINPUT111), .Z(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G124), .A2(n888), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n859), .B(KEYINPUT44), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT112), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G112), .A2(n890), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G100), .A2(n884), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G136), .A2(n885), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U967 ( .A(n867), .B(G160), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G130), .A2(n888), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G118), .A2(n890), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U972 ( .A1(n884), .A2(G106), .ZN(n872) );
  XOR2_X1 U973 ( .A(KEYINPUT113), .B(n872), .Z(n874) );
  NAND2_X1 U974 ( .A1(n885), .A2(G142), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(n918), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n900) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n882) );
  XNOR2_X1 U981 ( .A(G162), .B(KEYINPUT48), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(n883), .B(KEYINPUT116), .Z(n897) );
  NAND2_X1 U984 ( .A1(G103), .A2(n884), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n895) );
  NAND2_X1 U987 ( .A1(n888), .A2(G127), .ZN(n889) );
  XOR2_X1 U988 ( .A(KEYINPUT115), .B(n889), .Z(n892) );
  NAND2_X1 U989 ( .A1(G115), .A2(n890), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n930) );
  XNOR2_X1 U993 ( .A(n930), .B(KEYINPUT114), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U995 ( .A(G164), .B(n898), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n992), .B(n904), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(G171), .B(n905), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1002 ( .A(G286), .B(n908), .Z(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1004 ( .A(KEYINPUT110), .B(n910), .Z(G319) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n913) );
  AND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n915), .A2(G319), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1012 ( .A(G2084), .B(G160), .Z(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n924) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n922), .B(KEYINPUT51), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1021 ( .A(KEYINPUT118), .B(n929), .Z(n935) );
  XOR2_X1 U1022 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1025 ( .A(KEYINPUT50), .B(n933), .Z(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  NAND2_X1 U1029 ( .A1(n939), .A2(G29), .ZN(n1019) );
  XOR2_X1 U1030 ( .A(G25), .B(G1991), .Z(n940) );
  NAND2_X1 U1031 ( .A1(n940), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1032 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(G27), .B(n943), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1040 ( .A(KEYINPUT53), .B(n950), .Z(n953) );
  XOR2_X1 U1041 ( .A(KEYINPUT54), .B(G34), .Z(n951) );
  XNOR2_X1 U1042 ( .A(G2084), .B(n951), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1044 ( .A(KEYINPUT119), .B(G2090), .Z(n954) );
  XNOR2_X1 U1045 ( .A(G35), .B(n954), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(n957), .B(KEYINPUT120), .ZN(n958) );
  NOR2_X1 U1048 ( .A1(G29), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(KEYINPUT55), .B(n959), .ZN(n960) );
  NAND2_X1 U1050 ( .A1(n960), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1051 ( .A(G1966), .B(G21), .Z(n968) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G1976), .B(G23), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1055 ( .A(KEYINPUT126), .B(n963), .Z(n965) );
  XNOR2_X1 U1056 ( .A(G1986), .B(G24), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n981) );
  XOR2_X1 U1060 ( .A(G1961), .B(G5), .Z(n979) );
  XNOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n969), .B(G4), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(G1956), .B(G20), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1067 ( .A(KEYINPUT125), .B(G1341), .Z(n974) );
  XNOR2_X1 U1068 ( .A(G19), .B(n974), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n977), .B(KEYINPUT60), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT61), .B(n982), .Z(n983) );
  NOR2_X1 U1074 ( .A1(G16), .A2(n983), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT127), .B(n984), .ZN(n1015) );
  XOR2_X1 U1076 ( .A(G168), .B(G1966), .Z(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT121), .B(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n988), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G171), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1348), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1010) );
  INV_X1 U1086 ( .A(G1971), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(G166), .A2(n997), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT122), .B(n1002), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1003), .B(G1956), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1096 ( .A(G16), .B(KEYINPUT56), .Z(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(KEYINPUT124), .B(n1013), .Z(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1100 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

