

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764;

  INV_X2 U367 ( .A(G953), .ZN(n747) );
  NOR2_X1 U368 ( .A1(G953), .A2(G237), .ZN(n494) );
  XNOR2_X1 U369 ( .A(G137), .B(G128), .ZN(n383) );
  XNOR2_X1 U370 ( .A(n378), .B(KEYINPUT33), .ZN(n511) );
  INV_X1 U371 ( .A(G128), .ZN(n410) );
  NAND2_X1 U372 ( .A1(n399), .A2(n611), .ZN(n640) );
  NAND2_X2 U373 ( .A1(n366), .A2(n363), .ZN(n553) );
  NOR2_X2 U374 ( .A1(n356), .A2(n355), .ZN(n615) );
  AND2_X2 U375 ( .A1(n683), .A2(n358), .ZN(n355) );
  XNOR2_X2 U376 ( .A(n641), .B(n491), .ZN(n677) );
  AND2_X1 U377 ( .A1(n504), .A2(n481), .ZN(n386) );
  XNOR2_X1 U378 ( .A(n557), .B(KEYINPUT39), .ZN(n385) );
  AND2_X1 U379 ( .A1(n630), .A2(n581), .ZN(n373) );
  OR2_X1 U380 ( .A1(n585), .A2(n635), .ZN(n630) );
  XNOR2_X1 U381 ( .A(n354), .B(KEYINPUT73), .ZN(n556) );
  NAND2_X1 U382 ( .A1(n552), .A2(n551), .ZN(n354) );
  AND2_X1 U383 ( .A1(n368), .A2(n367), .ZN(n366) );
  XNOR2_X2 U384 ( .A(n347), .B(G469), .ZN(n377) );
  NOR2_X1 U385 ( .A1(n677), .A2(G902), .ZN(n347) );
  AND2_X1 U386 ( .A1(n673), .A2(n669), .ZN(n348) );
  NAND2_X1 U387 ( .A1(n517), .A2(n516), .ZN(n408) );
  XNOR2_X2 U388 ( .A(n359), .B(n601), .ZN(n399) );
  XNOR2_X1 U389 ( .A(n590), .B(n427), .ZN(n578) );
  NAND2_X1 U390 ( .A1(n553), .A2(n697), .ZN(n590) );
  NOR2_X1 U391 ( .A1(n362), .A2(n537), .ZN(n538) );
  AND2_X1 U392 ( .A1(n387), .A2(n351), .ZN(n362) );
  AND2_X1 U393 ( .A1(n370), .A2(n586), .ZN(n587) );
  INV_X1 U394 ( .A(n424), .ZN(n365) );
  NAND2_X1 U395 ( .A1(n424), .A2(n422), .ZN(n367) );
  XNOR2_X1 U396 ( .A(n507), .B(KEYINPUT66), .ZN(n525) );
  XNOR2_X1 U397 ( .A(G125), .B(G140), .ZN(n458) );
  XNOR2_X1 U398 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n457) );
  XNOR2_X1 U399 ( .A(G131), .B(G137), .ZN(n482) );
  XNOR2_X1 U400 ( .A(n464), .B(KEYINPUT99), .ZN(n699) );
  XNOR2_X1 U401 ( .A(n384), .B(n383), .ZN(n382) );
  XNOR2_X1 U402 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n384) );
  XNOR2_X1 U403 ( .A(n381), .B(G110), .ZN(n380) );
  XNOR2_X1 U404 ( .A(G119), .B(KEYINPUT91), .ZN(n381) );
  AND2_X1 U405 ( .A1(n569), .A2(n568), .ZN(n579) );
  NOR2_X2 U406 ( .A1(n578), .A2(n434), .ZN(n435) );
  INV_X1 U407 ( .A(KEYINPUT83), .ZN(n407) );
  NAND2_X1 U408 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U409 ( .A(KEYINPUT44), .ZN(n406) );
  NAND2_X1 U410 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U411 ( .A(G237), .ZN(n423) );
  XNOR2_X1 U412 ( .A(G116), .B(G101), .ZN(n417) );
  INV_X1 U413 ( .A(KEYINPUT2), .ZN(n358) );
  XNOR2_X1 U414 ( .A(G146), .B(KEYINPUT4), .ZN(n483) );
  XNOR2_X1 U415 ( .A(n402), .B(n401), .ZN(n400) );
  INV_X1 U416 ( .A(KEYINPUT17), .ZN(n401) );
  NAND2_X1 U417 ( .A1(n747), .A2(G224), .ZN(n402) );
  AND2_X1 U418 ( .A1(n598), .A2(n745), .ZN(n599) );
  INV_X1 U419 ( .A(n525), .ZN(n508) );
  NAND2_X1 U420 ( .A1(n365), .A2(n612), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n377), .B(n492), .ZN(n509) );
  INV_X1 U422 ( .A(KEYINPUT1), .ZN(n492) );
  OR2_X1 U423 ( .A1(n654), .A2(G902), .ZN(n398) );
  XNOR2_X1 U424 ( .A(KEYINPUT87), .B(G110), .ZN(n414) );
  NAND2_X1 U425 ( .A1(n640), .A2(n358), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n562), .B(KEYINPUT41), .ZN(n726) );
  XNOR2_X1 U427 ( .A(n515), .B(KEYINPUT35), .ZN(n539) );
  NAND2_X1 U428 ( .A1(n579), .A2(n374), .ZN(n585) );
  BUF_X1 U429 ( .A(n509), .Z(n493) );
  BUF_X1 U430 ( .A(n506), .Z(n708) );
  XNOR2_X1 U431 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U432 ( .A(n382), .B(n380), .ZN(n472) );
  XNOR2_X1 U433 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U434 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U435 ( .A(n661), .B(n662), .ZN(n663) );
  BUF_X1 U436 ( .A(n539), .Z(n671) );
  XNOR2_X1 U437 ( .A(n369), .B(n388), .ZN(n387) );
  INV_X1 U438 ( .A(KEYINPUT31), .ZN(n388) );
  NOR2_X1 U439 ( .A1(n717), .A2(n520), .ZN(n369) );
  INV_X1 U440 ( .A(G146), .ZN(n741) );
  AND2_X1 U441 ( .A1(n628), .A2(n665), .ZN(G66) );
  AND2_X1 U442 ( .A1(n611), .A2(KEYINPUT2), .ZN(n350) );
  NAND2_X1 U443 ( .A1(n638), .A2(n635), .ZN(n351) );
  AND2_X1 U444 ( .A1(n505), .A2(n481), .ZN(n352) );
  XNOR2_X1 U445 ( .A(G902), .B(KEYINPUT15), .ZN(n612) );
  NAND2_X1 U446 ( .A1(KEYINPUT83), .A2(KEYINPUT44), .ZN(n353) );
  NAND2_X1 U447 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X2 U448 ( .A(n526), .B(KEYINPUT93), .ZN(n552) );
  NAND2_X1 U449 ( .A1(n357), .A2(n422), .ZN(n356) );
  XNOR2_X1 U450 ( .A(n542), .B(n541), .ZN(n683) );
  NAND2_X1 U451 ( .A1(n600), .A2(n599), .ZN(n359) );
  XNOR2_X2 U452 ( .A(n360), .B(n560), .ZN(n670) );
  NAND2_X1 U453 ( .A1(n385), .A2(n591), .ZN(n360) );
  NAND2_X1 U454 ( .A1(n584), .A2(n371), .ZN(n370) );
  AND2_X2 U455 ( .A1(n673), .A2(n669), .ZN(n517) );
  NAND2_X1 U456 ( .A1(n361), .A2(n403), .ZN(n396) );
  INV_X1 U457 ( .A(n408), .ZN(n361) );
  XNOR2_X2 U458 ( .A(n435), .B(KEYINPUT0), .ZN(n510) );
  OR2_X2 U459 ( .A1(n525), .A2(n377), .ZN(n526) );
  NAND2_X1 U460 ( .A1(n404), .A2(n393), .ZN(n392) );
  OR2_X1 U461 ( .A1(n660), .A2(n364), .ZN(n363) );
  NAND2_X1 U462 ( .A1(n660), .A2(n424), .ZN(n368) );
  INV_X1 U463 ( .A(n742), .ZN(n372) );
  INV_X1 U464 ( .A(n578), .ZN(n374) );
  XNOR2_X2 U465 ( .A(n375), .B(KEYINPUT32), .ZN(n669) );
  NAND2_X1 U466 ( .A1(n535), .A2(n386), .ZN(n375) );
  XNOR2_X2 U467 ( .A(n376), .B(KEYINPUT100), .ZN(n673) );
  NAND2_X1 U468 ( .A1(n535), .A2(n352), .ZN(n376) );
  XNOR2_X2 U469 ( .A(n469), .B(n468), .ZN(n535) );
  XNOR2_X1 U470 ( .A(n377), .B(KEYINPUT103), .ZN(n569) );
  INV_X1 U471 ( .A(n511), .ZN(n727) );
  NAND2_X1 U472 ( .A1(n379), .A2(n593), .ZN(n378) );
  INV_X1 U473 ( .A(n518), .ZN(n379) );
  NAND2_X1 U474 ( .A1(n385), .A2(n529), .ZN(n603) );
  INV_X1 U475 ( .A(n556), .ZN(n577) );
  AND2_X1 U476 ( .A1(n387), .A2(n591), .ZN(n639) );
  AND2_X1 U477 ( .A1(n387), .A2(n529), .ZN(n637) );
  XNOR2_X1 U478 ( .A(n348), .B(KEYINPUT84), .ZN(n390) );
  NAND2_X1 U479 ( .A1(n391), .A2(n389), .ZN(n542) );
  NAND2_X1 U480 ( .A1(n540), .A2(n390), .ZN(n389) );
  NAND2_X1 U481 ( .A1(n394), .A2(n392), .ZN(n391) );
  OR2_X1 U482 ( .A1(n538), .A2(KEYINPUT83), .ZN(n393) );
  NAND2_X1 U483 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U484 ( .A1(n408), .A2(n353), .ZN(n395) );
  XNOR2_X2 U485 ( .A(n444), .B(G134), .ZN(n485) );
  XNOR2_X2 U486 ( .A(n397), .B(n410), .ZN(n444) );
  XNOR2_X2 U487 ( .A(G143), .B(KEYINPUT64), .ZN(n397) );
  NAND2_X1 U488 ( .A1(n714), .A2(n697), .ZN(n543) );
  XNOR2_X2 U489 ( .A(n398), .B(n501), .ZN(n714) );
  XNOR2_X1 U490 ( .A(n500), .B(n499), .ZN(n654) );
  NAND2_X1 U491 ( .A1(n399), .A2(n350), .ZN(n613) );
  XNOR2_X1 U492 ( .A(n444), .B(n400), .ZN(n413) );
  NAND2_X1 U493 ( .A1(n538), .A2(n407), .ZN(n403) );
  NAND2_X1 U494 ( .A1(n538), .A2(n405), .ZN(n404) );
  XNOR2_X2 U495 ( .A(n500), .B(KEYINPUT90), .ZN(n641) );
  AND2_X1 U496 ( .A1(n699), .A2(n707), .ZN(n409) );
  INV_X1 U497 ( .A(KEYINPUT46), .ZN(n573) );
  INV_X1 U498 ( .A(G122), .ZN(n440) );
  NAND2_X1 U499 ( .A1(n511), .A2(n510), .ZN(n513) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(G125), .B(KEYINPUT18), .ZN(n411) );
  XNOR2_X1 U502 ( .A(n483), .B(n411), .ZN(n412) );
  XNOR2_X1 U503 ( .A(n413), .B(n412), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n414), .B(G107), .ZN(n754) );
  XNOR2_X1 U505 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n415) );
  XNOR2_X1 U506 ( .A(n754), .B(n415), .ZN(n490) );
  XNOR2_X1 U507 ( .A(n416), .B(n490), .ZN(n421) );
  XNOR2_X1 U508 ( .A(n417), .B(G119), .ZN(n419) );
  XNOR2_X1 U509 ( .A(G113), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U510 ( .A(n419), .B(n418), .ZN(n498) );
  XNOR2_X1 U511 ( .A(G122), .B(G104), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n450), .B(KEYINPUT16), .ZN(n420) );
  XNOR2_X1 U513 ( .A(n498), .B(n420), .ZN(n755) );
  XNOR2_X1 U514 ( .A(n421), .B(n755), .ZN(n660) );
  INV_X1 U515 ( .A(n612), .ZN(n422) );
  INV_X1 U516 ( .A(G902), .ZN(n475) );
  NAND2_X1 U517 ( .A1(n423), .A2(n475), .ZN(n425) );
  AND2_X1 U518 ( .A1(n425), .A2(G210), .ZN(n424) );
  NAND2_X1 U519 ( .A1(n425), .A2(G214), .ZN(n426) );
  XNOR2_X1 U520 ( .A(n426), .B(KEYINPUT88), .ZN(n697) );
  INV_X1 U521 ( .A(KEYINPUT19), .ZN(n427) );
  NAND2_X1 U522 ( .A1(G234), .A2(G237), .ZN(n428) );
  XNOR2_X1 U523 ( .A(n428), .B(KEYINPUT14), .ZN(n431) );
  NAND2_X1 U524 ( .A1(G952), .A2(n431), .ZN(n725) );
  NOR2_X1 U525 ( .A1(G953), .A2(n725), .ZN(n429) );
  XNOR2_X1 U526 ( .A(n429), .B(KEYINPUT89), .ZN(n546) );
  AND2_X1 U527 ( .A1(G953), .A2(G902), .ZN(n430) );
  NAND2_X1 U528 ( .A1(n431), .A2(n430), .ZN(n544) );
  INV_X1 U529 ( .A(n544), .ZN(n432) );
  INV_X1 U530 ( .A(G898), .ZN(n756) );
  NAND2_X1 U531 ( .A1(n432), .A2(n756), .ZN(n433) );
  AND2_X1 U532 ( .A1(n546), .A2(n433), .ZN(n434) );
  XOR2_X1 U533 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n439) );
  NAND2_X1 U534 ( .A1(n747), .A2(G234), .ZN(n437) );
  INV_X1 U535 ( .A(KEYINPUT8), .ZN(n436) );
  XNOR2_X1 U536 ( .A(n437), .B(n436), .ZN(n470) );
  NAND2_X1 U537 ( .A1(G217), .A2(n470), .ZN(n438) );
  XNOR2_X1 U538 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U539 ( .A(G116), .B(G107), .ZN(n441) );
  XNOR2_X1 U540 ( .A(n445), .B(n485), .ZN(n650) );
  NAND2_X1 U541 ( .A1(n650), .A2(n475), .ZN(n447) );
  INV_X1 U542 ( .A(G478), .ZN(n446) );
  XNOR2_X1 U543 ( .A(n447), .B(n446), .ZN(n522) );
  NAND2_X1 U544 ( .A1(n494), .A2(G214), .ZN(n449) );
  XNOR2_X1 U545 ( .A(G143), .B(G131), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n449), .B(n448), .ZN(n452) );
  INV_X1 U547 ( .A(n450), .ZN(n451) );
  XNOR2_X1 U548 ( .A(n452), .B(n451), .ZN(n456) );
  XNOR2_X1 U549 ( .A(G113), .B(KEYINPUT12), .ZN(n454) );
  XNOR2_X1 U550 ( .A(KEYINPUT96), .B(KEYINPUT11), .ZN(n453) );
  XNOR2_X1 U551 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U552 ( .A(n456), .B(n455), .ZN(n459) );
  XNOR2_X1 U553 ( .A(n458), .B(n457), .ZN(n642) );
  XNOR2_X1 U554 ( .A(n642), .B(n741), .ZN(n473) );
  XNOR2_X1 U555 ( .A(n459), .B(n473), .ZN(n619) );
  OR2_X1 U556 ( .A1(n619), .A2(G902), .ZN(n463) );
  XNOR2_X1 U557 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n461) );
  XNOR2_X1 U558 ( .A(G475), .B(KEYINPUT97), .ZN(n460) );
  XNOR2_X1 U559 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U560 ( .A(n463), .B(n462), .ZN(n521) );
  INV_X1 U561 ( .A(n521), .ZN(n523) );
  NAND2_X1 U562 ( .A1(n522), .A2(n523), .ZN(n464) );
  NAND2_X1 U563 ( .A1(G234), .A2(n612), .ZN(n465) );
  XNOR2_X1 U564 ( .A(KEYINPUT20), .B(n465), .ZN(n476) );
  AND2_X1 U565 ( .A1(n476), .A2(G221), .ZN(n467) );
  XNOR2_X1 U566 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n467), .B(n466), .ZN(n707) );
  NAND2_X1 U568 ( .A1(n510), .A2(n409), .ZN(n469) );
  XNOR2_X1 U569 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n468) );
  NAND2_X1 U570 ( .A1(n470), .A2(G221), .ZN(n471) );
  XNOR2_X1 U571 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n474), .B(n473), .ZN(n627) );
  NAND2_X1 U573 ( .A1(n627), .A2(n475), .ZN(n480) );
  XOR2_X1 U574 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n478) );
  NAND2_X1 U575 ( .A1(n476), .A2(G217), .ZN(n477) );
  XNOR2_X1 U576 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X2 U577 ( .A(n480), .B(n479), .ZN(n506) );
  INV_X1 U578 ( .A(n708), .ZN(n481) );
  XNOR2_X1 U579 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X2 U580 ( .A(n485), .B(n484), .ZN(n500) );
  NAND2_X1 U581 ( .A1(n747), .A2(G227), .ZN(n486) );
  XNOR2_X1 U582 ( .A(n486), .B(G140), .ZN(n488) );
  XNOR2_X1 U583 ( .A(G101), .B(G104), .ZN(n487) );
  XNOR2_X1 U584 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U585 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U586 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n496) );
  NAND2_X1 U587 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U589 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U590 ( .A(G472), .B(KEYINPUT70), .ZN(n501) );
  INV_X1 U591 ( .A(KEYINPUT6), .ZN(n502) );
  XNOR2_X1 U592 ( .A(n714), .B(n502), .ZN(n593) );
  XNOR2_X1 U593 ( .A(n593), .B(KEYINPUT75), .ZN(n503) );
  AND2_X1 U594 ( .A1(n493), .A2(n503), .ZN(n504) );
  INV_X1 U595 ( .A(n493), .ZN(n711) );
  INV_X1 U596 ( .A(n714), .ZN(n528) );
  AND2_X1 U597 ( .A1(n711), .A2(n528), .ZN(n505) );
  NAND2_X1 U598 ( .A1(n506), .A2(n707), .ZN(n507) );
  NAND2_X1 U599 ( .A1(n509), .A2(n508), .ZN(n518) );
  INV_X1 U600 ( .A(KEYINPUT34), .ZN(n512) );
  XNOR2_X1 U601 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U602 ( .A(n522), .ZN(n524) );
  AND2_X1 U603 ( .A1(n524), .A2(n521), .ZN(n575) );
  NAND2_X1 U604 ( .A1(n514), .A2(n575), .ZN(n515) );
  INV_X1 U605 ( .A(n539), .ZN(n516) );
  NOR2_X1 U606 ( .A1(n518), .A2(n528), .ZN(n519) );
  XNOR2_X1 U607 ( .A(n519), .B(KEYINPUT95), .ZN(n717) );
  INV_X1 U608 ( .A(n510), .ZN(n520) );
  AND2_X1 U609 ( .A1(n522), .A2(n521), .ZN(n591) );
  INV_X1 U610 ( .A(n591), .ZN(n638) );
  AND2_X1 U611 ( .A1(n524), .A2(n523), .ZN(n529) );
  INV_X1 U612 ( .A(n529), .ZN(n635) );
  NAND2_X1 U613 ( .A1(n510), .A2(n552), .ZN(n531) );
  NAND2_X1 U614 ( .A1(n591), .A2(n528), .ZN(n527) );
  NOR2_X1 U615 ( .A1(n531), .A2(n527), .ZN(n737) );
  NAND2_X1 U616 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U617 ( .A1(n531), .A2(n530), .ZN(n739) );
  NOR2_X1 U618 ( .A1(n737), .A2(n739), .ZN(n536) );
  INV_X1 U619 ( .A(n593), .ZN(n532) );
  NAND2_X1 U620 ( .A1(n532), .A2(n708), .ZN(n533) );
  NOR2_X1 U621 ( .A1(n493), .A2(n533), .ZN(n534) );
  NAND2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n633) );
  NAND2_X1 U623 ( .A1(n536), .A2(n633), .ZN(n537) );
  NOR2_X1 U624 ( .A1(n671), .A2(KEYINPUT44), .ZN(n540) );
  XOR2_X1 U625 ( .A(KEYINPUT80), .B(KEYINPUT45), .Z(n541) );
  XNOR2_X1 U626 ( .A(n543), .B(KEYINPUT30), .ZN(n550) );
  XOR2_X1 U627 ( .A(KEYINPUT101), .B(n544), .Z(n545) );
  OR2_X1 U628 ( .A1(G900), .A2(n545), .ZN(n547) );
  NAND2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U630 ( .A(KEYINPUT76), .ZN(n548) );
  XNOR2_X1 U631 ( .A(n549), .B(n548), .ZN(n563) );
  NOR2_X1 U632 ( .A1(n550), .A2(n563), .ZN(n551) );
  BUF_X1 U633 ( .A(n553), .Z(n554) );
  XNOR2_X1 U634 ( .A(n554), .B(KEYINPUT38), .ZN(n700) );
  INV_X1 U635 ( .A(n700), .ZN(n555) );
  XNOR2_X1 U636 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n559) );
  INV_X1 U637 ( .A(KEYINPUT106), .ZN(n558) );
  XNOR2_X1 U638 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U639 ( .A1(n699), .A2(n697), .ZN(n561) );
  OR2_X1 U640 ( .A1(n561), .A2(n700), .ZN(n562) );
  NOR2_X1 U641 ( .A1(n506), .A2(n563), .ZN(n564) );
  AND2_X1 U642 ( .A1(n707), .A2(n564), .ZN(n592) );
  NAND2_X1 U643 ( .A1(n714), .A2(n592), .ZN(n567) );
  XNOR2_X1 U644 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n565) );
  XNOR2_X1 U645 ( .A(n565), .B(KEYINPUT28), .ZN(n566) );
  XNOR2_X1 U646 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U647 ( .A1(n726), .A2(n579), .ZN(n571) );
  INV_X1 U648 ( .A(KEYINPUT42), .ZN(n570) );
  XNOR2_X1 U649 ( .A(n571), .B(n570), .ZN(n764) );
  INV_X1 U650 ( .A(n764), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n670), .A2(n572), .ZN(n574) );
  XNOR2_X1 U652 ( .A(n574), .B(n573), .ZN(n600) );
  NAND2_X1 U653 ( .A1(n575), .A2(n554), .ZN(n576) );
  OR2_X1 U654 ( .A1(n577), .A2(n576), .ZN(n632) );
  NOR2_X1 U655 ( .A1(n585), .A2(n638), .ZN(n742) );
  INV_X1 U656 ( .A(KEYINPUT47), .ZN(n580) );
  AND2_X1 U657 ( .A1(n580), .A2(KEYINPUT78), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n585), .A2(KEYINPUT78), .ZN(n583) );
  AND2_X1 U659 ( .A1(n351), .A2(KEYINPUT47), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U661 ( .A1(n585), .A2(KEYINPUT78), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n632), .A2(n587), .ZN(n589) );
  INV_X1 U663 ( .A(KEYINPUT72), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n589), .B(n588), .ZN(n598) );
  AND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n604) );
  NOR2_X1 U667 ( .A1(n590), .A2(n604), .ZN(n596) );
  XNOR2_X1 U668 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n596), .B(n595), .ZN(n597) );
  OR2_X1 U670 ( .A1(n711), .A2(n597), .ZN(n745) );
  INV_X1 U671 ( .A(KEYINPUT48), .ZN(n601) );
  INV_X1 U672 ( .A(KEYINPUT108), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n603), .B(n602), .ZN(n762) );
  INV_X1 U674 ( .A(n604), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n697), .A2(n605), .ZN(n606) );
  OR2_X1 U676 ( .A1(n493), .A2(n606), .ZN(n608) );
  XNOR2_X1 U677 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n608), .B(n607), .ZN(n610) );
  INV_X1 U679 ( .A(n554), .ZN(n609) );
  AND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n634) );
  NOR2_X1 U681 ( .A1(n762), .A2(n634), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT81), .ZN(n614) );
  INV_X1 U683 ( .A(n683), .ZN(n748) );
  NAND2_X1 U684 ( .A1(n614), .A2(n748), .ZN(n692) );
  NAND2_X1 U685 ( .A1(n615), .A2(n692), .ZN(n616) );
  XNOR2_X2 U686 ( .A(n616), .B(KEYINPUT65), .ZN(n674) );
  NAND2_X1 U687 ( .A1(n674), .A2(G475), .ZN(n621) );
  XNOR2_X1 U688 ( .A(KEYINPUT86), .B(KEYINPUT122), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT59), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U691 ( .A(G952), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n622), .A2(G953), .ZN(n665) );
  NAND2_X1 U693 ( .A1(n623), .A2(n665), .ZN(n625) );
  INV_X1 U694 ( .A(KEYINPUT60), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(G60) );
  NAND2_X1 U696 ( .A1(n674), .A2(G217), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(n628) );
  INV_X1 U698 ( .A(n665), .ZN(n680) );
  XOR2_X1 U699 ( .A(G128), .B(KEYINPUT29), .Z(n629) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G30) );
  XOR2_X1 U701 ( .A(G143), .B(KEYINPUT111), .Z(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(G45) );
  XNOR2_X1 U703 ( .A(n633), .B(G101), .ZN(G3) );
  XOR2_X1 U704 ( .A(G140), .B(n634), .Z(G42) );
  XNOR2_X1 U705 ( .A(G116), .B(KEYINPUT113), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(G18) );
  XOR2_X1 U707 ( .A(G113), .B(n639), .Z(G15) );
  XNOR2_X1 U708 ( .A(n642), .B(KEYINPUT125), .ZN(n643) );
  XNOR2_X1 U709 ( .A(n641), .B(n643), .ZN(n645) );
  XNOR2_X1 U710 ( .A(n640), .B(n645), .ZN(n644) );
  NAND2_X1 U711 ( .A1(n644), .A2(n747), .ZN(n649) );
  XNOR2_X1 U712 ( .A(G227), .B(n645), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n646), .A2(G900), .ZN(n647) );
  NAND2_X1 U714 ( .A1(n647), .A2(G953), .ZN(n648) );
  NAND2_X1 U715 ( .A1(n649), .A2(n648), .ZN(G72) );
  NAND2_X1 U716 ( .A1(n674), .A2(G478), .ZN(n651) );
  XOR2_X1 U717 ( .A(n651), .B(n650), .Z(n652) );
  NOR2_X1 U718 ( .A1(n652), .A2(n680), .ZN(G63) );
  NAND2_X1 U719 ( .A1(n674), .A2(G472), .ZN(n656) );
  XNOR2_X1 U720 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n657), .A2(n665), .ZN(n659) );
  XNOR2_X1 U723 ( .A(KEYINPUT110), .B(KEYINPUT63), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n659), .B(n658), .ZN(G57) );
  NAND2_X1 U725 ( .A1(n674), .A2(G210), .ZN(n664) );
  BUF_X1 U726 ( .A(n660), .Z(n661) );
  XNOR2_X1 U727 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n664), .B(n663), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n667) );
  XNOR2_X1 U731 ( .A(n668), .B(n667), .ZN(G51) );
  XNOR2_X1 U732 ( .A(n669), .B(G119), .ZN(G21) );
  XNOR2_X1 U733 ( .A(n670), .B(G131), .ZN(G33) );
  XNOR2_X1 U734 ( .A(G122), .B(KEYINPUT126), .ZN(n672) );
  XOR2_X1 U735 ( .A(n672), .B(n671), .Z(G24) );
  XNOR2_X1 U736 ( .A(n673), .B(G110), .ZN(G12) );
  NAND2_X1 U737 ( .A1(n674), .A2(G469), .ZN(n679) );
  XNOR2_X1 U738 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n675) );
  XNOR2_X1 U739 ( .A(n675), .B(KEYINPUT58), .ZN(n676) );
  XNOR2_X1 U740 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n679), .B(n678), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(G54) );
  INV_X1 U743 ( .A(n640), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n682), .A2(KEYINPUT79), .ZN(n685) );
  BUF_X1 U745 ( .A(n683), .Z(n684) );
  NOR2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U747 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n687) );
  NOR2_X1 U748 ( .A1(n686), .A2(n687), .ZN(n691) );
  INV_X1 U749 ( .A(n687), .ZN(n688) );
  NAND2_X1 U750 ( .A1(n640), .A2(n688), .ZN(n689) );
  AND2_X1 U751 ( .A1(n689), .A2(KEYINPUT79), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n733) );
  XNOR2_X1 U754 ( .A(n700), .B(KEYINPUT117), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n699), .A2(n694), .ZN(n696) );
  INV_X1 U756 ( .A(n697), .ZN(n695) );
  NAND2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n704) );
  NAND2_X1 U758 ( .A1(n697), .A2(KEYINPUT117), .ZN(n698) );
  NAND2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U760 ( .A1(n351), .A2(n555), .ZN(n701) );
  NAND2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U763 ( .A1(n727), .A2(n705), .ZN(n706) );
  XNOR2_X1 U764 ( .A(n706), .B(KEYINPUT118), .ZN(n722) );
  NOR2_X1 U765 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U766 ( .A(n709), .B(KEYINPUT49), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n710), .B(KEYINPUT116), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n711), .A2(n525), .ZN(n712) );
  XOR2_X1 U769 ( .A(KEYINPUT50), .B(n712), .Z(n713) );
  NOR2_X1 U770 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U771 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U772 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(n719), .Z(n720) );
  NAND2_X1 U774 ( .A1(n720), .A2(n726), .ZN(n721) );
  NAND2_X1 U775 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U776 ( .A(KEYINPUT52), .B(n723), .Z(n724) );
  NOR2_X1 U777 ( .A1(n725), .A2(n724), .ZN(n730) );
  INV_X1 U778 ( .A(n726), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U781 ( .A(KEYINPUT119), .B(n731), .Z(n732) );
  NAND2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n734), .B(KEYINPUT120), .ZN(n735) );
  NOR2_X1 U784 ( .A1(n735), .A2(G953), .ZN(n736) );
  XNOR2_X1 U785 ( .A(n736), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U786 ( .A(G104), .B(n737), .Z(G6) );
  XNOR2_X1 U787 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U789 ( .A(G107), .B(n740), .ZN(G9) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U791 ( .A(KEYINPUT112), .B(n743), .ZN(G48) );
  XOR2_X1 U792 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U794 ( .A(G125), .B(n746), .ZN(G27) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(n753) );
  NAND2_X1 U796 ( .A1(G953), .A2(G224), .ZN(n749) );
  XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n749), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G898), .ZN(n751) );
  XOR2_X1 U799 ( .A(KEYINPUT123), .B(n751), .Z(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n760) );
  XNOR2_X1 U801 ( .A(n755), .B(n754), .ZN(n758) );
  NAND2_X1 U802 ( .A1(n756), .A2(G953), .ZN(n757) );
  AND2_X1 U803 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U804 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U805 ( .A(KEYINPUT124), .B(n761), .ZN(G69) );
  XNOR2_X1 U806 ( .A(G134), .B(KEYINPUT115), .ZN(n763) );
  XNOR2_X1 U807 ( .A(n763), .B(n762), .ZN(G36) );
  XOR2_X1 U808 ( .A(n764), .B(G137), .Z(G39) );
endmodule

