//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT92), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n204), .B(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT92), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT15), .B(new_n203), .C1(new_n209), .C2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n207), .B2(new_n208), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT93), .B1(new_n215), .B2(G50gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n217), .B(new_n203), .Z(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G1gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G1gat), .B2(new_n220), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(G8gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT94), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n219), .B(KEYINPUT17), .ZN(new_n227));
  INV_X1    g026(.A(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT18), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n226), .A2(new_n229), .A3(KEYINPUT18), .A4(new_n230), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n219), .A2(new_n224), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT95), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n225), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT95), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n235), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n230), .B(KEYINPUT13), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n233), .B(new_n234), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT11), .B(G169gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  INV_X1    g047(.A(KEYINPUT96), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n233), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n243), .A2(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n202), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n243), .A2(new_n250), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT97), .A3(new_n251), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  XNOR2_X1  g058(.A(G15gat), .B(G43gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G71gat), .B(G99gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G227gat), .ZN(new_n264));
  INV_X1    g063(.A(G233gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT23), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT24), .A3(new_n269), .ZN(new_n275));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n271), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n271), .A2(KEYINPUT64), .A3(new_n275), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n267), .A2(KEYINPUT23), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n277), .A2(KEYINPUT25), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(KEYINPUT25), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n271), .A2(new_n275), .A3(new_n279), .A4(new_n276), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n273), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n273), .B1(new_n289), .B2(KEYINPUT65), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n286), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n267), .A2(KEYINPUT26), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n292), .A2(new_n269), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n305), .A3(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n301), .ZN(new_n308));
  OR2_X1    g107(.A1(G127gat), .A2(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT66), .B(G127gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n296), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n284), .B2(new_n296), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n266), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n319), .B(new_n266), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT33), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n263), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n316), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n314), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n319), .B1(new_n326), .B2(new_n266), .ZN(new_n327));
  INV_X1    g126(.A(new_n320), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT32), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n266), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n325), .A2(new_n330), .A3(new_n314), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT34), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT34), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n325), .A2(new_n333), .A3(new_n330), .A4(new_n314), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n334), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(KEYINPUT32), .B2(new_n321), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n324), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n335), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n321), .A3(KEYINPUT32), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n323), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n343), .B(KEYINPUT36), .Z(new_n344));
  AND2_X1   g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n284), .A2(new_n296), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT69), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G197gat), .B(G204gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT70), .ZN(new_n356));
  XOR2_X1   g155(.A(G211gat), .B(G218gat), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n355), .B2(new_n356), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n350), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT71), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n345), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n346), .A2(KEYINPUT72), .A3(new_n345), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n348), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n372), .B2(new_n366), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  INV_X1    g173(.A(G64gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G92gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT30), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n372), .A2(new_n366), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n378), .B1(new_n382), .B2(new_n367), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n373), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n385), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT0), .B(G57gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G85gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n307), .A2(new_n312), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT73), .ZN(new_n395));
  AND2_X1   g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G155gat), .ZN(new_n399));
  INV_X1    g198(.A(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT73), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(KEYINPUT2), .ZN(new_n405));
  INV_X1    g204(.A(G148gat), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n406), .A2(G141gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(G141gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT74), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT75), .B(G162gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G155gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT2), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n407), .A2(new_n408), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n402), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n394), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n404), .A2(new_n412), .A3(new_n409), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n412), .B1(new_n404), .B2(new_n409), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n394), .B(new_n420), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n393), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n431), .B2(new_n313), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n430), .A2(new_n393), .A3(KEYINPUT79), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(KEYINPUT76), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n424), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT80), .A3(new_n393), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n428), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT81), .B1(new_n441), .B2(KEYINPUT5), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n443), .B(new_n444), .C1(new_n438), .C2(new_n440), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT3), .B1(new_n421), .B2(new_n425), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n452));
  AND4_X1   g251(.A1(new_n393), .A2(new_n448), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n430), .A2(new_n393), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n439), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n442), .A2(new_n445), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n448), .A2(new_n393), .A3(new_n451), .A4(new_n452), .ZN(new_n461));
  INV_X1    g260(.A(new_n433), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT79), .B1(new_n430), .B2(new_n393), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n456), .A2(new_n454), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n440), .A2(KEYINPUT5), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT82), .A4(new_n467), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n392), .B1(new_n460), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT80), .B1(new_n436), .B2(new_n393), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n427), .B(new_n313), .C1(new_n435), .C2(new_n424), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n439), .B1(new_n477), .B2(new_n434), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n443), .B1(new_n478), .B2(new_n444), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n441), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n461), .A2(new_n439), .A3(new_n457), .A4(new_n455), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n470), .A2(new_n471), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n391), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n473), .A2(new_n474), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT6), .B(new_n392), .C1(new_n460), .C2(new_n472), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n387), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n360), .A2(new_n361), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n347), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n363), .A2(new_n488), .A3(new_n347), .A4(new_n359), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n436), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT29), .B1(new_n431), .B2(new_n450), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n365), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n494), .A2(new_n496), .A3(G228gat), .A4(G233gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n357), .A2(KEYINPUT83), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n353), .A2(new_n498), .A3(new_n354), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n357), .A2(KEYINPUT83), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n347), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n355), .A2(new_n500), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n450), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n430), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n365), .B2(new_n495), .ZN(new_n505));
  INV_X1    g304(.A(G228gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n265), .ZN(new_n507));
  INV_X1    g306(.A(G22gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n497), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G78gat), .B(G106gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT31), .ZN(new_n511));
  INV_X1    g310(.A(G50gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT85), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n507), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G22gat), .ZN(new_n518));
  AOI211_X1 g317(.A(new_n508), .B(new_n513), .C1(new_n497), .C2(new_n507), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n509), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n509), .A2(new_n515), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT86), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n344), .B1(new_n487), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n486), .A2(KEYINPUT88), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n391), .B1(new_n482), .B2(new_n483), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT6), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n482), .A2(new_n391), .A3(new_n483), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n526), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n525), .A2(new_n528), .B1(new_n530), .B2(new_n474), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT38), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n385), .A2(KEYINPUT37), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n379), .B1(new_n373), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n372), .A2(new_n366), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(KEYINPUT37), .C1(new_n366), .C2(new_n349), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n532), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n383), .B1(new_n536), .B2(new_n537), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n531), .A2(new_n539), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n520), .A2(new_n521), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n461), .A2(new_n466), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n440), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT39), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(new_n392), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(KEYINPUT39), .C1(new_n440), .C2(new_n438), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT40), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n387), .A2(new_n473), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n551), .A2(new_n552), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n555), .A2(KEYINPUT40), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n547), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n524), .B1(new_n546), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n547), .A2(new_n559), .A3(new_n343), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n487), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n340), .A2(new_n323), .A3(new_n341), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n323), .B1(new_n340), .B2(new_n341), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n339), .A2(KEYINPUT90), .A3(new_n342), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n522), .B1(new_n386), .B2(new_n384), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n525), .A2(new_n528), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n485), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n561), .B1(new_n570), .B2(KEYINPUT35), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n259), .B1(new_n558), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n569), .A2(new_n485), .A3(new_n544), .A4(new_n545), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n557), .B1(new_n573), .B2(new_n538), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n343), .B(KEYINPUT36), .ZN(new_n575));
  INV_X1    g374(.A(new_n487), .ZN(new_n576));
  INV_X1    g375(.A(new_n523), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n485), .A2(new_n486), .ZN(new_n580));
  INV_X1    g379(.A(new_n387), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n560), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n569), .A2(new_n485), .ZN(new_n583));
  INV_X1    g382(.A(new_n567), .ZN(new_n584));
  INV_X1    g383(.A(new_n568), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n586), .B2(new_n559), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n258), .B1(new_n572), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G71gat), .B(G78gat), .Z(new_n590));
  AOI21_X1  g389(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n375), .A2(G57gat), .ZN(new_n593));
  INV_X1    g392(.A(G57gat), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n594), .A2(KEYINPUT99), .A3(G64gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT99), .B1(new_n594), .B2(G64gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(G64gat), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n599), .A2(new_n593), .A3(KEYINPUT98), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT98), .B1(new_n599), .B2(new_n593), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n600), .A2(new_n601), .A3(new_n591), .ZN(new_n602));
  INV_X1    g401(.A(new_n590), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n224), .B1(new_n605), .B2(KEYINPUT21), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G183gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G127gat), .B(G155gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n612), .B(new_n616), .Z(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(G85gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n618), .B1(new_n619), .B2(new_n377), .ZN(new_n620));
  NAND2_X1  g419(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n619), .B2(new_n377), .ZN(new_n622));
  NAND4_X1  g421(.A1(KEYINPUT101), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G99gat), .B(G106gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n227), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n219), .A2(new_n626), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G134gat), .B(G162gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT102), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  XOR2_X1   g436(.A(new_n633), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n604), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n626), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n626), .B1(new_n605), .B2(KEYINPUT103), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n627), .A2(new_n604), .A3(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT104), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(KEYINPUT105), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n643), .B1(new_n640), .B2(new_n626), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n646), .B1(new_n654), .B2(new_n642), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n655), .B2(new_n650), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n654), .A2(new_n651), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  INV_X1    g458(.A(G176gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G204gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n651), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n657), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n617), .A2(new_n638), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n589), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n580), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g473(.A1(new_n670), .A2(new_n581), .ZN(new_n675));
  INV_X1    g474(.A(G8gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n221), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n221), .A2(new_n676), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT42), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1325gat));
  AND3_X1   g483(.A1(new_n671), .A2(G15gat), .A3(new_n575), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n671), .B2(new_n584), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n670), .A2(new_n523), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n688), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(new_n617), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n668), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n589), .A2(new_n638), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n207), .A4(new_n672), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n589), .A2(new_n672), .A3(new_n638), .A4(new_n693), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT45), .B1(new_n697), .B2(G29gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n638), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n572), .B2(new_n588), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n579), .A2(new_n587), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n705), .B2(new_n638), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n255), .A2(new_n251), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n693), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n704), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(KEYINPUT108), .A3(new_n672), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n587), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT91), .B1(new_n579), .B2(new_n587), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n702), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n705), .A2(new_n638), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n701), .ZN(new_n715));
  INV_X1    g514(.A(new_n708), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n713), .A2(new_n672), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n710), .A2(G29gat), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n699), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n699), .A2(new_n720), .A3(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n694), .A2(new_n208), .A3(new_n387), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n727));
  INV_X1    g526(.A(new_n709), .ZN(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n728), .B2(new_n581), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n728), .B2(new_n344), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n709), .A2(KEYINPUT110), .A3(new_n575), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(G43gat), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n694), .A2(new_n215), .A3(new_n584), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(KEYINPUT47), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  INV_X1    g537(.A(new_n736), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n215), .B1(new_n709), .B2(new_n575), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(G1330gat));
  AOI21_X1  g541(.A(new_n512), .B1(new_n709), .B2(new_n577), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n589), .A2(new_n512), .A3(new_n638), .A4(new_n693), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n523), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n713), .A2(new_n547), .A3(new_n715), .A4(new_n716), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G50gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n693), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n258), .B(new_n750), .C1(new_n572), .C2(new_n588), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n751), .A2(new_n512), .A3(new_n577), .A4(new_n638), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n744), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT111), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n713), .A2(new_n577), .A3(new_n715), .A4(new_n716), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n744), .A3(new_n752), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  INV_X1    g557(.A(new_n745), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n759), .A2(new_n577), .B1(new_n748), .B2(G50gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n757), .B(new_n758), .C1(new_n760), .C2(new_n744), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n754), .A2(new_n761), .ZN(G1331gat));
  INV_X1    g561(.A(new_n668), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n707), .B(new_n763), .C1(new_n579), .C2(new_n587), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n617), .A2(new_n638), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n580), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT112), .B(G57gat), .Z(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1332gat));
  NOR2_X1   g568(.A1(new_n766), .A2(new_n581), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  AND2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n770), .B2(new_n771), .ZN(G1333gat));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n766), .A2(new_n775), .A3(new_n344), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n764), .A2(new_n584), .A3(new_n765), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g578(.A1(new_n766), .A2(new_n523), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g580(.A1(new_n692), .A2(new_n707), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n704), .A2(new_n706), .A3(new_n763), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(G85gat), .A3(new_n672), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n714), .B2(new_n783), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n705), .A2(new_n787), .A3(new_n638), .A4(new_n782), .ZN(new_n788));
  AND4_X1   g587(.A1(new_n672), .A2(new_n786), .A3(new_n668), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n789), .B2(G85gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1336gat));
  NAND3_X1  g591(.A1(new_n784), .A2(G92gat), .A3(new_n387), .ZN(new_n793));
  AND4_X1   g592(.A1(new_n387), .A2(new_n786), .A3(new_n668), .A4(new_n788), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n795), .B(new_n796), .ZN(G1337gat));
  NAND2_X1  g596(.A1(new_n784), .A2(new_n575), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n798), .A2(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(G99gat), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n567), .A2(G99gat), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n668), .A3(new_n788), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1338gat));
  INV_X1    g603(.A(G106gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n784), .B2(new_n577), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n786), .A2(new_n547), .A3(new_n668), .A4(new_n788), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(G106gat), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT53), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n807), .B2(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n784), .A2(new_n547), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n810), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n805), .B1(new_n784), .B2(new_n547), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n812), .A3(KEYINPUT115), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n809), .B1(new_n816), .B2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT105), .B1(new_n648), .B2(new_n651), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n655), .A2(new_n653), .A3(new_n650), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n820), .B(new_n663), .C1(new_n823), .C2(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT54), .B1(new_n652), .B2(new_n656), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT117), .B1(new_n825), .B2(new_n666), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n648), .A2(KEYINPUT116), .A3(new_n651), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(new_n648), .B2(new_n651), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n665), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n824), .A2(new_n826), .A3(KEYINPUT55), .A4(new_n829), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n707), .A3(new_n667), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n241), .A2(new_n242), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n226), .A2(new_n229), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(G229gat), .A3(G233gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n247), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n243), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n248), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n668), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n638), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n832), .A2(new_n667), .A3(new_n833), .A4(new_n840), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n700), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n617), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n669), .A2(new_n255), .A3(new_n251), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(KEYINPUT118), .A3(new_n846), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n523), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n580), .A2(new_n387), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n584), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n258), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n857));
  AND4_X1   g656(.A1(new_n672), .A2(new_n851), .A3(new_n342), .A4(new_n339), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n585), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n707), .A2(new_n299), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT120), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n856), .A2(new_n857), .B1(new_n859), .B2(new_n861), .ZN(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n854), .B2(new_n763), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n858), .A2(new_n297), .A3(new_n585), .A4(new_n668), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n311), .A3(new_n617), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n858), .A2(new_n585), .A3(new_n692), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n311), .B2(new_n871), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n638), .A2(new_n310), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT56), .B1(new_n859), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT122), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n859), .A2(KEYINPUT56), .A3(new_n873), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n854), .B2(new_n700), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n878), .B(KEYINPUT56), .C1(new_n859), .C2(new_n873), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n879), .ZN(G1343gat));
  NAND3_X1  g679(.A1(new_n849), .A2(new_n547), .A3(new_n850), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n853), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n575), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n257), .A2(new_n667), .A3(new_n832), .A4(new_n833), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n638), .B1(new_n888), .B2(new_n841), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n617), .B1(new_n889), .B2(new_n844), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n846), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n577), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894), .B2(new_n258), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n882), .A2(new_n886), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n258), .A2(G141gat), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  INV_X1    g699(.A(new_n894), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n707), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(G141gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n903), .B2(new_n896), .ZN(G1344gat));
  NAND2_X1  g703(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n669), .A2(new_n258), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n577), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n905), .A2(new_n668), .A3(new_n886), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n881), .A2(KEYINPUT57), .B1(new_n907), .B2(new_n577), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(KEYINPUT124), .A3(new_n668), .A4(new_n886), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(G148gat), .A3(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n406), .C1(new_n901), .C2(new_n668), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n668), .A2(new_n406), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n916), .A2(new_n917), .B1(new_n897), .B2(new_n918), .ZN(G1345gat));
  NOR3_X1   g718(.A1(new_n894), .A2(new_n399), .A3(new_n617), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n882), .A2(new_n692), .A3(new_n886), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n399), .B2(new_n921), .ZN(G1346gat));
  NOR2_X1   g721(.A1(new_n897), .A2(new_n700), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n415), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n901), .A2(new_n415), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n638), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n672), .A2(new_n581), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n852), .A2(new_n584), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n258), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n849), .A2(new_n850), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n547), .A3(new_n343), .ZN(new_n933));
  INV_X1    g732(.A(G169gat), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n707), .A4(new_n927), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT125), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n931), .A3(new_n936), .ZN(G1348gat));
  NOR3_X1   g736(.A1(new_n928), .A2(new_n660), .A3(new_n763), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n933), .A2(new_n927), .ZN(new_n939));
  AOI21_X1  g738(.A(G176gat), .B1(new_n939), .B2(new_n668), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n933), .A2(new_n285), .A3(new_n692), .A4(new_n927), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n851), .A2(new_n523), .A3(new_n584), .ZN(new_n943));
  INV_X1    g742(.A(new_n927), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n943), .A2(new_n617), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n945), .B2(new_n272), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n939), .A2(new_n273), .A3(new_n638), .ZN(new_n948));
  OAI21_X1  g747(.A(G190gat), .B1(new_n928), .B2(new_n700), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n944), .A2(new_n575), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n881), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(G197gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(new_n707), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT127), .ZN(new_n958));
  INV_X1    g757(.A(new_n912), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(new_n258), .A3(new_n954), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n958), .B1(new_n956), .B2(new_n960), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n955), .A2(new_n662), .A3(new_n668), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n959), .A2(new_n763), .A3(new_n954), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n963), .B(new_n964), .C1(new_n965), .C2(new_n662), .ZN(G1353gat));
  INV_X1    g765(.A(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n955), .A2(new_n967), .A3(new_n692), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n912), .A2(new_n692), .A3(new_n953), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  INV_X1    g771(.A(G218gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n973), .A3(new_n638), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n959), .A2(new_n700), .A3(new_n954), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n973), .ZN(G1355gat));
endmodule


