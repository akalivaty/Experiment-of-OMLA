//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939;
  INV_X1    g000(.A(G226gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n209), .B1(new_n216), .B2(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(KEYINPUT65), .B2(new_n216), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI211_X1 g019(.A(new_n219), .B(new_n209), .C1(new_n215), .C2(new_n210), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT28), .A3(new_n214), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT27), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G183gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(new_n214), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT66), .A4(new_n214), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n227), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n236), .ZN(new_n238));
  AOI211_X1 g037(.A(KEYINPUT68), .B(new_n238), .C1(new_n233), .C2(new_n234), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n226), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT69), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(new_n226), .C1(new_n237), .C2(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n205), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n246));
  INV_X1    g045(.A(new_n207), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n224), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  AOI211_X1 g049(.A(KEYINPUT70), .B(new_n248), .C1(new_n241), .C2(new_n243), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n204), .B(new_n223), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n225), .B2(new_n214), .ZN(new_n253));
  AND4_X1   g052(.A1(KEYINPUT66), .A2(new_n228), .A3(new_n230), .A4(new_n214), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n236), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n235), .A2(new_n227), .A3(new_n236), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n242), .B1(new_n258), .B2(new_n226), .ZN(new_n259));
  INV_X1    g058(.A(new_n226), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT69), .B(new_n260), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n249), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n223), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n204), .A2(KEYINPUT29), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT77), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n273), .B2(KEYINPUT76), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(KEYINPUT76), .B2(new_n273), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT78), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT78), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n282), .A3(new_n279), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n223), .A2(new_n204), .A3(new_n262), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n248), .B1(new_n241), .B2(new_n243), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n224), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n222), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n264), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n284), .B(new_n287), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(new_n293), .A3(new_n297), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT30), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G155gat), .B(G162gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G141gat), .B(G148gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n304), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT2), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G113gat), .B(G120gat), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n316), .B2(KEYINPUT1), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n321));
  NAND4_X1  g120(.A1(new_n318), .A2(new_n315), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n312), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n317), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n311), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT81), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n324), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n325), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  OR3_X1    g139(.A1(new_n339), .A2(KEYINPUT39), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT0), .ZN(new_n343));
  XNOR2_X1  g142(.A(G57gat), .B(G85gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NOR2_X1   g144(.A1(new_n339), .A2(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n329), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n323), .ZN(new_n348));
  INV_X1    g147(.A(new_n340), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT39), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n341), .B(new_n345), .C1(new_n346), .C2(new_n350), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n351), .A2(KEYINPUT40), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(KEYINPUT40), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n294), .A2(KEYINPUT30), .A3(new_n298), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT86), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT5), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n348), .B2(new_n349), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n331), .B2(new_n333), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n340), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n334), .A2(new_n357), .A3(new_n340), .A4(new_n338), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n345), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n356), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT86), .B(new_n345), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n301), .A2(new_n354), .A3(new_n355), .A4(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT37), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n291), .A2(new_n204), .B1(new_n264), .B2(new_n263), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n293), .B(new_n370), .C1(new_n371), .C2(new_n284), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n286), .A2(KEYINPUT87), .A3(new_n370), .A4(new_n293), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT38), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n298), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n287), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n223), .B1(new_n250), .B2(new_n251), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n264), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n370), .B1(new_n381), .B2(new_n285), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n266), .A2(new_n284), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n364), .A2(new_n365), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n364), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT6), .B1(new_n389), .B2(new_n345), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n368), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n300), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n370), .B1(new_n286), .B2(new_n293), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(new_n297), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n377), .B1(new_n376), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n369), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n277), .B1(new_n275), .B2(new_n273), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(new_n335), .B1(new_n330), .B2(new_n328), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n312), .B2(new_n335), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n281), .B2(new_n283), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n400), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n405), .B(KEYINPUT84), .ZN(new_n408));
  OAI211_X1 g207(.A(G228gat), .B(G233gat), .C1(new_n285), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT83), .B1(new_n280), .B2(new_n402), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n280), .A2(KEYINPUT83), .A3(new_n402), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n312), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n399), .B(new_n407), .C1(new_n409), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT85), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n407), .B1(new_n409), .B2(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G22gat), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT31), .B(G50gat), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT82), .ZN(new_n419));
  XOR2_X1   g218(.A(G78gat), .B(G106gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AND4_X1   g220(.A1(new_n414), .A2(new_n415), .A3(new_n417), .A4(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n415), .A2(new_n421), .B1(new_n417), .B2(new_n414), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n398), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n388), .B1(new_n386), .B2(new_n390), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n301), .B2(new_n355), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n422), .A2(new_n423), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT36), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n380), .A2(new_n326), .ZN(new_n433));
  INV_X1    g232(.A(G227gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n203), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n325), .B(new_n223), .C1(new_n250), .C2(new_n251), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT73), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n444), .A2(KEYINPUT74), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(KEYINPUT74), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT33), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(KEYINPUT32), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT34), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n436), .ZN(new_n453));
  INV_X1    g252(.A(new_n435), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT34), .B(new_n435), .C1(new_n433), .C2(new_n436), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n446), .A3(new_n450), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n432), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n455), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n453), .A2(new_n452), .A3(new_n454), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n446), .A2(new_n450), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT75), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(new_n460), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(KEYINPUT75), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n461), .B1(new_n467), .B2(new_n432), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n427), .A2(new_n424), .A3(new_n459), .A4(new_n460), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n301), .A2(new_n355), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n391), .A2(KEYINPUT35), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n471), .A2(new_n424), .A3(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n457), .A2(new_n446), .A3(new_n450), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n474), .A2(new_n464), .A3(KEYINPUT75), .ZN(new_n475));
  INV_X1    g274(.A(new_n465), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n431), .A2(new_n468), .B1(new_n470), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479));
  OR2_X1    g278(.A1(G43gat), .A2(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G43gat), .A2(G50gat), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT89), .B(G50gat), .Z(new_n483));
  OAI211_X1 g282(.A(new_n479), .B(new_n481), .C1(new_n483), .C2(G43gat), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT14), .B(G29gat), .Z(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(G36gat), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n482), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(G1gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498));
  AOI21_X1  g297(.A(G8gat), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT92), .A3(KEYINPUT16), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT16), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(G1gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n496), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n497), .B(new_n505), .C1(new_n498), .C2(G8gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT17), .B1(new_n489), .B2(new_n490), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n509), .B(KEYINPUT94), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n491), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT95), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT88), .B(G197gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT11), .B(G169gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT12), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n513), .B(new_n491), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n512), .B(KEYINPUT13), .Z(new_n526));
  AOI22_X1  g325(.A1(new_n515), .A2(new_n516), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n511), .A2(KEYINPUT18), .A3(new_n512), .A4(new_n514), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n527), .B(new_n528), .C1(new_n517), .C2(new_n523), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n478), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT96), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT98), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(KEYINPUT98), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n513), .B1(new_n542), .B2(KEYINPUT21), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT99), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n538), .B(KEYINPUT96), .Z(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n547));
  AND2_X1   g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G127gat), .B(G155gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT97), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n549), .B(new_n551), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n549), .B(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n544), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n555), .A3(new_n559), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n570), .B2(new_n571), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G99gat), .B(G106gat), .Z(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n495), .A2(new_n510), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT101), .Z(new_n583));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n581), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n586), .A2(new_n491), .B1(KEYINPUT41), .B2(new_n564), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n585), .B1(new_n583), .B2(new_n587), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n568), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n567), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G230gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n203), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n586), .A2(KEYINPUT10), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n540), .B2(new_n541), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n546), .A2(new_n581), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n538), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT10), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n600), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n605), .ZN(new_n609));
  INV_X1    g408(.A(new_n600), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n598), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n602), .B2(new_n606), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n613), .B(new_n597), .C1(new_n610), .C2(new_n609), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(KEYINPUT102), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n616), .B(new_n598), .C1(new_n608), .C2(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n563), .A2(new_n594), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n563), .A2(new_n594), .A3(KEYINPUT103), .A4(new_n618), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n533), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n426), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n500), .ZN(G1324gat));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(new_n471), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT16), .B(G8gat), .Z(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(G8gat), .B1(new_n624), .B2(new_n471), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  MUX2_X1   g432(.A(new_n631), .B(new_n633), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g433(.A(G15gat), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n624), .A2(new_n635), .A3(new_n468), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n628), .A2(new_n467), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT104), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(new_n640), .A3(new_n635), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(G1326gat));
  NOR2_X1   g441(.A1(new_n624), .A2(new_n424), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT43), .B(G22gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n477), .A2(new_n470), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n432), .B1(new_n475), .B2(new_n476), .ZN(new_n647));
  INV_X1    g446(.A(new_n461), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n429), .B1(new_n398), .B2(new_n424), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n532), .ZN(new_n652));
  INV_X1    g451(.A(new_n618), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n563), .A2(new_n594), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(G29gat), .A3(new_n625), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT45), .Z(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n478), .B2(new_n594), .ZN(new_n659));
  INV_X1    g458(.A(new_n594), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(KEYINPUT44), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n561), .A2(KEYINPUT105), .A3(new_n562), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT105), .B1(new_n561), .B2(new_n562), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n532), .A3(new_n653), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT106), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668), .B2(new_n625), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n657), .A2(new_n669), .ZN(G1328gat));
  OAI21_X1  g469(.A(G36gat), .B1(new_n668), .B2(new_n471), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n655), .A2(G36gat), .A3(new_n471), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT46), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n667), .A3(new_n649), .A4(new_n661), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G43gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n467), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n655), .A2(G43gat), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1330gat));
  NAND4_X1  g480(.A1(new_n659), .A2(new_n667), .A3(new_n428), .A4(new_n661), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n483), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n533), .A2(KEYINPUT107), .A3(new_n654), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n655), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n424), .A2(new_n483), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT108), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1331gat));
  INV_X1    g491(.A(new_n563), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n693), .A2(new_n660), .A3(new_n652), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n653), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(new_n651), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n426), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n651), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n471), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  AND2_X1   g502(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n702), .B2(new_n703), .ZN(G1333gat));
  INV_X1    g505(.A(G71gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n701), .B2(new_n677), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n468), .A2(new_n707), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT110), .B1(new_n698), .B2(new_n709), .ZN(new_n710));
  AND4_X1   g509(.A1(KEYINPUT110), .A2(new_n697), .A3(new_n651), .A4(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT50), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n714), .B(new_n708), .C1(new_n710), .C2(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1334gat));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n424), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT111), .B(G78gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n563), .A2(new_n652), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n653), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT112), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n662), .A2(new_n426), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n651), .A2(new_n660), .A3(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n720), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n725), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n651), .A2(new_n660), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n651), .A2(KEYINPUT113), .A3(new_n660), .A4(new_n728), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n726), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n653), .A2(new_n570), .A3(new_n426), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT114), .ZN(new_n736));
  OAI22_X1  g535(.A1(new_n723), .A2(new_n570), .B1(new_n734), .B2(new_n736), .ZN(G1336gat));
  NAND4_X1  g536(.A1(new_n659), .A2(new_n629), .A3(new_n661), .A4(new_n722), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT52), .B1(new_n738), .B2(G92gat), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n471), .A2(G92gat), .A3(new_n618), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n392), .B1(new_n376), .B2(new_n384), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n297), .B(new_n395), .C1(new_n374), .C2(new_n375), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n377), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n428), .B1(new_n745), .B2(new_n369), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n648), .B(new_n647), .C1(new_n746), .C2(new_n429), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n594), .B(new_n727), .C1(new_n747), .C2(new_n646), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT116), .B1(new_n748), .B2(KEYINPUT51), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n750), .A3(new_n725), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n729), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n740), .B(KEYINPUT115), .Z(new_n753));
  AOI22_X1  g552(.A1(new_n752), .A2(new_n753), .B1(G92gat), .B2(new_n738), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n742), .B1(new_n754), .B2(new_n755), .ZN(G1337gat));
  NOR3_X1   g555(.A1(new_n677), .A2(G99gat), .A3(new_n618), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n659), .A2(new_n649), .A3(new_n661), .A4(new_n722), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n733), .A2(new_n757), .B1(new_n758), .B2(G99gat), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1338gat));
  NAND4_X1  g560(.A1(new_n659), .A2(new_n428), .A3(new_n661), .A4(new_n722), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT53), .B1(new_n762), .B2(G106gat), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n424), .A2(G106gat), .A3(new_n618), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n730), .A2(new_n729), .B1(new_n724), .B2(new_n725), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n732), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n767), .B2(KEYINPUT118), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n733), .A2(KEYINPUT118), .A3(new_n764), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n752), .A2(new_n764), .B1(G106gat), .B2(new_n762), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(G1339gat));
  AND4_X1   g571(.A1(new_n532), .A2(new_n563), .A3(new_n594), .A4(new_n618), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n603), .A2(new_n607), .A3(new_n600), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n776), .A2(new_n613), .A3(KEYINPUT54), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n598), .B1(new_n613), .B2(KEYINPUT54), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n597), .B1(new_n608), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(new_n613), .A3(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT55), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n614), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n525), .A2(new_n526), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n512), .B1(new_n511), .B2(new_n514), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n522), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT119), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n527), .A2(new_n523), .A3(new_n528), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n522), .C1(new_n786), .C2(new_n787), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n785), .A2(new_n591), .A3(new_n593), .A4(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n532), .A2(new_n784), .B1(new_n618), .B2(new_n793), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n660), .B1(KEYINPUT120), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799));
  OAI221_X1 g598(.A(new_n799), .B1(new_n618), .B2(new_n793), .C1(new_n532), .C2(new_n784), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n796), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n774), .B1(new_n801), .B2(new_n665), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n677), .A2(new_n428), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n629), .A2(new_n625), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(G113gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n532), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n797), .A2(KEYINPUT120), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n594), .A3(new_n800), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n665), .B1(new_n810), .B2(new_n795), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n625), .B1(new_n812), .B2(new_n774), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n466), .A2(new_n428), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n652), .A3(new_n471), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n808), .B1(new_n807), .B2(new_n816), .ZN(G1340gat));
  INV_X1    g616(.A(G120gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n806), .A2(new_n818), .A3(new_n618), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n471), .A3(new_n653), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n818), .B2(new_n820), .ZN(G1341gat));
  INV_X1    g620(.A(new_n665), .ZN(new_n822));
  OAI21_X1  g621(.A(G127gat), .B1(new_n806), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n815), .A2(new_n471), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n693), .A2(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(G1342gat));
  NAND2_X1  g625(.A1(new_n660), .A2(new_n471), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(G134gat), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n802), .A2(new_n426), .A3(new_n814), .A4(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n802), .A2(new_n660), .A3(new_n805), .A4(new_n803), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT121), .B1(new_n832), .B2(G134gat), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n832), .A2(KEYINPUT121), .A3(G134gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n831), .B(KEYINPUT122), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n649), .A2(new_n424), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n813), .A2(new_n471), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(G141gat), .A3(new_n532), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(KEYINPUT58), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n428), .C1(new_n811), .C2(new_n773), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n468), .A2(new_n805), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n797), .A2(new_n594), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n563), .B1(new_n848), .B2(new_n795), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n428), .B1(new_n849), .B2(new_n773), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G141gat), .B1(new_n852), .B2(new_n532), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n843), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n845), .A2(new_n851), .A3(KEYINPUT123), .A4(new_n847), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n652), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n842), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(G1344gat));
  OR3_X1    g660(.A1(new_n841), .A2(G148gat), .A3(new_n618), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G148gat), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n856), .A2(new_n857), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n653), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n802), .A2(new_n428), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n621), .A2(new_n532), .A3(new_n622), .ZN(new_n868));
  INV_X1    g667(.A(new_n849), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n424), .A2(KEYINPUT57), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n867), .A2(KEYINPUT57), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n653), .A3(new_n847), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n863), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n862), .B1(new_n866), .B2(new_n874), .ZN(G1345gat));
  NOR3_X1   g674(.A1(new_n841), .A2(KEYINPUT124), .A3(new_n693), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(G155gat), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT124), .B1(new_n841), .B2(new_n693), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n822), .A2(new_n308), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n877), .A2(new_n878), .B1(new_n865), .B2(new_n879), .ZN(G1346gat));
  NOR2_X1   g679(.A1(new_n827), .A2(G162gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n813), .A2(new_n840), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n865), .A2(new_n660), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n309), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n471), .A2(new_n426), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n804), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886), .B2(new_n532), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n811), .A2(new_n773), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n426), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n466), .A2(new_n471), .A3(new_n428), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n532), .A2(G169gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR4_X1   g696(.A1(new_n894), .A2(KEYINPUT126), .A3(G169gat), .A4(new_n532), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n887), .B1(new_n897), .B2(new_n898), .ZN(G1348gat));
  OAI21_X1  g698(.A(G176gat), .B1(new_n886), .B2(new_n618), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n618), .A2(G176gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n894), .B2(new_n901), .ZN(G1349gat));
  OAI21_X1  g701(.A(G183gat), .B1(new_n886), .B2(new_n822), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n563), .A2(new_n225), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n894), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT60), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n903), .B(new_n907), .C1(new_n894), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n895), .A2(new_n214), .A3(new_n660), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n804), .A2(new_n660), .A3(new_n885), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(G190gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n911), .B2(G190gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G1351gat));
  AND3_X1   g714(.A1(new_n890), .A2(new_n629), .A3(new_n840), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n652), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n468), .A2(new_n885), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n872), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n652), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n923), .A3(new_n653), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n872), .A2(new_n653), .A3(new_n919), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G204gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n916), .A2(new_n269), .A3(new_n563), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n872), .A2(new_n563), .A3(new_n919), .ZN(new_n932));
  AND4_X1   g731(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n269), .B1(KEYINPUT127), .B2(new_n934), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n932), .A2(new_n935), .B1(new_n931), .B2(KEYINPUT63), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n930), .B1(new_n933), .B2(new_n936), .ZN(G1354gat));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n270), .A3(new_n660), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n920), .A2(new_n660), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n270), .ZN(G1355gat));
endmodule


