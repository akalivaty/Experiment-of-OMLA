//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  AOI21_X1  g003(.A(G131), .B1(new_n188), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n190), .A3(KEYINPUT65), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(new_n192), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n191), .A2(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(G131), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(new_n203), .A3(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT64), .B1(new_n205), .B2(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G146), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n206), .A2(new_n209), .A3(G128), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G143), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n202), .A2(new_n204), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n211), .A2(KEYINPUT1), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n188), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n222), .B2(new_n199), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n197), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G116), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n231), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT28), .B1(new_n218), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n218), .A2(KEYINPUT67), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n202), .A2(new_n240), .A3(new_n204), .A4(new_n217), .ZN(new_n241));
  INV_X1    g055(.A(new_n224), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n235), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(new_n241), .A3(new_n236), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n238), .B1(new_n246), .B2(KEYINPUT28), .ZN(new_n247));
  NOR2_X1   g061(.A1(G237), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G210), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n249), .B(KEYINPUT27), .Z(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XOR2_X1   g065(.A(new_n250), .B(new_n251), .Z(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(KEYINPUT29), .ZN(new_n253));
  AOI21_X1  g067(.A(G902), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n224), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n239), .A2(new_n241), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n235), .ZN(new_n258));
  INV_X1    g072(.A(new_n201), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n242), .B1(new_n259), .B2(new_n216), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n245), .ZN(new_n263));
  INV_X1    g077(.A(new_n252), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT29), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n235), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n245), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n237), .B(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT70), .A4(new_n252), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n245), .B2(new_n266), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n238), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT70), .B1(new_n275), .B2(new_n252), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n254), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G472), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n268), .A2(new_n270), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n262), .A2(new_n245), .A3(new_n252), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n280), .A2(new_n264), .B1(KEYINPUT31), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n262), .A2(new_n283), .A3(new_n245), .A4(new_n252), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n245), .A2(new_n252), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n283), .A4(new_n262), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n279), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n292), .ZN(new_n294));
  AOI211_X1 g108(.A(KEYINPUT32), .B(new_n294), .C1(new_n282), .C2(new_n290), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n278), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G125), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G140), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n301), .A3(KEYINPUT73), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(KEYINPUT16), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G146), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n208), .A3(new_n305), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n225), .B2(G128), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n225), .A2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G110), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT24), .B(G110), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n225), .B2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n219), .A2(KEYINPUT71), .A3(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n313), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n309), .B(new_n316), .C1(new_n317), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n317), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n315), .B2(G110), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n298), .A2(new_n301), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n208), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n307), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n327), .A3(new_n332), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G217), .ZN(new_n337));
  INV_X1    g151(.A(G902), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(G234), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G902), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n341), .A2(KEYINPUT75), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n343), .B2(KEYINPUT74), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n334), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(KEYINPUT74), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n339), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(KEYINPUT75), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT9), .B(G234), .ZN(new_n353));
  OAI21_X1  g167(.A(G221), .B1(new_n353), .B2(G902), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT76), .ZN(new_n355));
  INV_X1    g169(.A(G469), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n338), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n330), .A2(G227), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT77), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G140), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(G104), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n365), .A2(G104), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(G107), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(G104), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n363), .B(new_n367), .C1(new_n370), .C2(KEYINPUT3), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G104), .B2(new_n365), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(KEYINPUT80), .A3(G107), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G107), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n384));
  INV_X1    g198(.A(new_n221), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  INV_X1    g203(.A(new_n368), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n391), .B2(new_n366), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n392), .A2(new_n371), .A3(KEYINPUT4), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(G101), .C1(new_n391), .C2(new_n366), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n217), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n395), .A2(new_n217), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n392), .A2(new_n371), .A3(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n386), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n202), .A2(new_n204), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n363), .B1(new_n376), .B2(new_n380), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n389), .A2(new_n390), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n366), .B1(new_n405), .B2(new_n364), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n406), .B2(new_n363), .ZN(new_n407));
  AND4_X1   g221(.A1(G128), .A2(new_n206), .A3(new_n209), .A4(new_n210), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n213), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G128), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT82), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT81), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n407), .A2(new_n418), .A3(KEYINPUT83), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT83), .B1(new_n407), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n384), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n402), .A2(new_n403), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n403), .B1(new_n402), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n362), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n407), .A2(new_n221), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n407), .A2(new_n418), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n407), .A2(new_n418), .A3(KEYINPUT83), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n426), .B1(new_n432), .B2(new_n403), .ZN(new_n433));
  INV_X1    g247(.A(new_n427), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n419), .B2(new_n420), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n436));
  NOR2_X1   g250(.A1(new_n259), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n422), .A3(new_n361), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n425), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n357), .B1(new_n441), .B2(new_n356), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n361), .ZN(new_n443));
  INV_X1    g257(.A(new_n403), .ZN(new_n444));
  INV_X1    g258(.A(new_n386), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n393), .A2(KEYINPUT79), .A3(new_n396), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n399), .B1(new_n398), .B2(new_n400), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT10), .B1(new_n430), .B2(new_n431), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT86), .B1(new_n422), .B2(new_n361), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT12), .B1(new_n435), .B2(new_n444), .ZN(new_n454));
  INV_X1    g268(.A(new_n437), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n432), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n422), .B(new_n453), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n362), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n453), .B1(new_n439), .B2(new_n422), .ZN(new_n459));
  OAI221_X1 g273(.A(G469), .B1(new_n451), .B2(new_n452), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n355), .B1(new_n442), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n230), .A2(KEYINPUT5), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g279(.A(G113), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n464), .A2(new_n467), .B1(new_n230), .B2(new_n232), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n371), .A3(new_n382), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n395), .A2(new_n235), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n393), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G122), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(new_n469), .C1(new_n393), .C2(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n216), .A2(G125), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(G125), .B2(new_n221), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n330), .A2(G224), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT87), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n480), .B(new_n482), .Z(new_n483));
  AND3_X1   g297(.A1(new_n476), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n469), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n407), .A2(KEYINPUT88), .A3(new_n468), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n487), .C1(new_n407), .C2(new_n468), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n472), .B(KEYINPUT8), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n482), .A2(KEYINPUT7), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n480), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n480), .A2(KEYINPUT89), .A3(new_n491), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT89), .B1(new_n480), .B2(new_n491), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n475), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n338), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT90), .B(new_n463), .C1(new_n484), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n476), .A2(new_n478), .A3(new_n483), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n493), .A2(new_n494), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n488), .A2(new_n489), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n475), .A4(new_n492), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n463), .A2(KEYINPUT90), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n498), .A2(new_n501), .A3(new_n338), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G214), .B1(G237), .B2(G902), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT93), .B1(new_n219), .B2(G143), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n205), .A3(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n219), .A2(G143), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n512), .A2(new_n188), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n188), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G116), .B(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n369), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT96), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n369), .A2(new_n517), .A3(KEYINPUT96), .ZN(new_n521));
  INV_X1    g335(.A(G122), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(new_n522), .B2(G116), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n227), .A3(G122), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n523), .B(new_n525), .C1(new_n227), .C2(G122), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n520), .A2(new_n521), .B1(G107), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n516), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(G107), .ZN(new_n530));
  INV_X1    g344(.A(new_n521), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT96), .B1(new_n369), .B2(new_n517), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n514), .A2(new_n515), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT97), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n514), .A2(KEYINPUT95), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n512), .A2(new_n188), .A3(new_n513), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n369), .A2(new_n517), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n537), .A2(new_n540), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n512), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT13), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n544), .B(new_n513), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n545), .ZN(new_n548));
  OAI21_X1  g362(.A(G134), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n536), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n353), .A2(new_n337), .A3(G953), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n529), .A2(new_n535), .B1(new_n542), .B2(new_n549), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n552), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(KEYINPUT98), .B(G902), .C1(new_n554), .C2(new_n556), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n508), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n248), .A2(G214), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n205), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n248), .A2(G143), .A3(G214), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G131), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT17), .ZN(new_n567));
  INV_X1    g381(.A(G131), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n568), .A3(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(KEYINPUT17), .A3(G131), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n307), .A2(new_n570), .A3(new_n308), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(KEYINPUT18), .A2(G131), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n563), .A2(new_n564), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n563), .B2(new_n564), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n299), .A2(G146), .A3(new_n302), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n326), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G113), .B(G122), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n374), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n572), .A2(new_n582), .A3(new_n579), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT92), .B(G475), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n585), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n306), .A2(G146), .B1(new_n566), .B2(new_n569), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT19), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n299), .B2(new_n302), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n325), .A2(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n208), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n590), .A2(new_n594), .B1(new_n578), .B2(new_n576), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n582), .B1(new_n595), .B2(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n566), .A2(new_n569), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n307), .A2(new_n597), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n579), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(G475), .A2(G902), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT20), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n583), .B1(new_n599), .B2(new_n600), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n585), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT20), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n603), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n588), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n555), .A2(new_n552), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n536), .A2(new_n550), .A3(new_n552), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n338), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n508), .B1(new_n614), .B2(KEYINPUT98), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n330), .A2(G952), .ZN(new_n617));
  INV_X1    g431(.A(G234), .ZN(new_n618));
  INV_X1    g432(.A(G237), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n338), .B(new_n330), .C1(G234), .C2(G237), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT21), .B(G898), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n561), .A2(new_n611), .A3(new_n616), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT99), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n614), .A2(KEYINPUT98), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n557), .A2(new_n558), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n615), .B1(new_n630), .B2(new_n508), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n611), .A4(new_n625), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n506), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n296), .A2(new_n352), .A3(new_n461), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n264), .B1(new_n238), .B2(new_n274), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n257), .A2(new_n261), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT31), .B1(new_n639), .B2(new_n286), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n289), .B2(new_n285), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n642), .B2(G902), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n294), .B1(new_n282), .B2(new_n290), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n645), .A3(new_n352), .ZN(new_n646));
  INV_X1    g460(.A(new_n461), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n637), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n462), .B1(new_n484), .B2(new_n496), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n498), .A2(new_n501), .A3(new_n338), .A4(new_n463), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n505), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n624), .ZN(new_n652));
  INV_X1    g466(.A(G472), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n291), .B2(new_n338), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n644), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n352), .A4(new_n461), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n554), .A2(new_n556), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n551), .A2(KEYINPUT101), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT33), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n554), .A2(new_n658), .A3(KEYINPUT33), .A4(new_n556), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n507), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n507), .A2(new_n338), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n614), .B2(G478), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n611), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n648), .A2(new_n652), .A3(new_n656), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NAND2_X1  g483(.A1(new_n648), .A2(new_n656), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n604), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n609), .B1(new_n608), .B2(new_n603), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n588), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n605), .A2(new_n675), .A3(new_n610), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n649), .A2(new_n505), .A3(new_n650), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n561), .A2(new_n616), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .A4(new_n625), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n670), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NOR2_X1   g497(.A1(new_n333), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n328), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n340), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n349), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n655), .A2(new_n634), .A3(new_n461), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  NAND3_X1  g505(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n621), .B1(new_n622), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n692), .A2(new_n631), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n422), .A2(new_n361), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n435), .A2(new_n444), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n697), .A2(new_n426), .B1(new_n435), .B2(new_n437), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n361), .B1(new_n450), .B2(new_n422), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n356), .B(new_n338), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n357), .ZN(new_n702));
  OAI22_X1  g516(.A1(new_n458), .A2(new_n459), .B1(new_n451), .B2(new_n452), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n356), .ZN(new_n704));
  INV_X1    g518(.A(new_n355), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n695), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n688), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n651), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n706), .A2(new_n296), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT104), .B(G128), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G30));
  OAI21_X1  g525(.A(new_n338), .B1(new_n246), .B2(new_n252), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n264), .B1(new_n262), .B2(new_n245), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n293), .B2(new_n295), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n504), .B(KEYINPUT38), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n611), .B1(new_n561), .B2(new_n616), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n707), .A2(new_n505), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n694), .B(KEYINPUT39), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n461), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  NAND2_X1  g541(.A1(new_n660), .A2(new_n661), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G478), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n674), .B1(new_n671), .B2(new_n672), .ZN(new_n730));
  INV_X1    g544(.A(new_n665), .ZN(new_n731));
  INV_X1    g545(.A(new_n694), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n355), .B(new_n733), .C1(new_n442), .C2(new_n460), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n296), .A2(new_n734), .A3(new_n708), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  OAI21_X1  g550(.A(KEYINPUT32), .B1(new_n642), .B2(new_n294), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n644), .A2(new_n279), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n351), .B1(new_n739), .B2(new_n278), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n338), .B1(new_n699), .B2(new_n700), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n701), .A3(new_n354), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n678), .A2(new_n666), .A3(new_n625), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR2_X1   g562(.A1(new_n680), .A2(new_n743), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NAND4_X1  g565(.A1(new_n742), .A2(new_n678), .A3(new_n701), .A4(new_n354), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n707), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n627), .A2(new_n633), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n296), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT105), .B(G119), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G21));
  OAI21_X1  g571(.A(new_n640), .B1(new_n247), .B2(new_n252), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(KEYINPUT106), .B(new_n640), .C1(new_n247), .C2(new_n252), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n290), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n654), .B1(new_n762), .B2(new_n292), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n652), .A2(new_n719), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n743), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n352), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NOR3_X1   g581(.A1(new_n752), .A2(new_n707), .A3(new_n733), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n763), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NAND3_X1  g584(.A1(new_n497), .A2(new_n505), .A3(new_n503), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n733), .A2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n704), .A2(new_n772), .A3(new_n354), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT42), .B1(new_n740), .B2(new_n773), .ZN(new_n774));
  AND4_X1   g588(.A1(KEYINPUT42), .A2(new_n773), .A3(new_n296), .A4(new_n352), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n568), .ZN(G33));
  AND2_X1   g591(.A1(new_n704), .A2(new_n354), .ZN(new_n778));
  INV_X1    g592(.A(new_n771), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n740), .A2(new_n695), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n356), .B1(new_n703), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n703), .A2(new_n782), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n783), .B2(KEYINPUT107), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n357), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n701), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n354), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n722), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n662), .A2(new_n665), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n611), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT43), .Z(new_n796));
  OAI211_X1 g610(.A(new_n796), .B(new_n688), .C1(new_n644), .C2(new_n654), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n771), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n191), .ZN(G39));
  OR2_X1    g616(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n739), .A2(new_n278), .A3(new_n351), .A4(new_n772), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT108), .B(G140), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G42));
  NAND3_X1  g624(.A1(new_n352), .A2(new_n705), .A3(new_n505), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n717), .A3(new_n795), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n742), .A2(new_n701), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n812), .A2(new_n716), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n635), .A2(new_n766), .A3(new_n689), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n296), .B(new_n352), .C1(new_n749), .C2(new_n745), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n755), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n506), .A2(new_n624), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n648), .A2(new_n656), .A3(new_n666), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n679), .A2(new_n611), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT109), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n648), .A2(new_n656), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n818), .A2(new_n820), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n773), .A2(new_n763), .A3(new_n688), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n688), .A2(new_n631), .A3(new_n732), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n692), .A3(new_n771), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n296), .A2(new_n461), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(new_n780), .C1(new_n774), .C2(new_n775), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n719), .A2(new_n678), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n688), .A3(new_n694), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n715), .A2(new_n778), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n735), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n708), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n739), .B2(new_n278), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n839), .A2(new_n706), .B1(new_n763), .B2(new_n768), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n709), .A2(new_n735), .A3(new_n836), .A4(new_n769), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT113), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n842), .A2(new_n843), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n833), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n709), .A2(new_n769), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n856));
  OAI211_X1 g670(.A(KEYINPUT52), .B(new_n837), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n847), .A2(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n847), .A2(KEYINPUT112), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n833), .A2(KEYINPUT110), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT110), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n826), .B2(new_n832), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n852), .B1(new_n864), .B2(KEYINPUT53), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n850), .A2(new_n869), .A3(new_n851), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n850), .B2(new_n851), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n866), .B1(new_n865), .B2(KEYINPUT54), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n743), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT118), .B1(new_n876), .B2(new_n779), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n743), .A2(new_n878), .A3(new_n771), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n620), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n796), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n881), .A2(new_n688), .A3(new_n763), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n796), .A2(new_n621), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n763), .A2(new_n352), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n717), .A2(new_n505), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n743), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT50), .Z(new_n888));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n880), .A2(new_n352), .A3(new_n716), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n794), .A2(new_n730), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n890), .A2(new_n889), .A3(new_n892), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n882), .B(new_n888), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n705), .B1(new_n813), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n896), .B2(new_n813), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n803), .A2(new_n804), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n885), .A2(new_n771), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT116), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n895), .A2(KEYINPUT51), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n881), .A2(new_n740), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT48), .Z(new_n908));
  INV_X1    g722(.A(new_n666), .ZN(new_n909));
  OAI221_X1 g723(.A(new_n617), .B1(new_n885), .B2(new_n752), .C1(new_n890), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n875), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n817), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NAND3_X1  g729(.A1(new_n872), .A2(G210), .A3(G902), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n476), .A2(new_n478), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(new_n483), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n917), .A2(new_n918), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n330), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n916), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n921), .B1(new_n930), .B2(KEYINPUT56), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(G51));
  XNOR2_X1  g746(.A(new_n872), .B(KEYINPUT54), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n357), .B(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n425), .A2(new_n440), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n850), .A2(new_n851), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT115), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n850), .A2(new_n869), .A3(new_n851), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n338), .B1(new_n941), .B2(new_n868), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n784), .A3(new_n786), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n928), .B1(new_n937), .B2(new_n943), .ZN(G54));
  NAND3_X1  g758(.A1(new_n942), .A2(KEYINPUT58), .A3(G475), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n945), .A2(new_n602), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n602), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n947), .A3(new_n928), .ZN(G60));
  INV_X1    g762(.A(new_n728), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n663), .B(KEYINPUT59), .Z(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n875), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n933), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n929), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n951), .A2(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n872), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n336), .B(KEYINPUT124), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n928), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n941), .B2(new_n868), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n686), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n962), .A2(new_n872), .A3(new_n686), .A4(new_n958), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(KEYINPUT61), .B(new_n961), .C1(new_n964), .C2(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G66));
  INV_X1    g784(.A(G224), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n623), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n826), .B(KEYINPUT125), .Z(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n919), .B1(G898), .B2(new_n330), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  NAND2_X1  g791(.A1(new_n260), .A2(new_n255), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n257), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n592), .A2(new_n593), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n856), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n982), .A2(new_n854), .B1(new_n839), .B2(new_n734), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n726), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  AOI21_X1  g799(.A(new_n801), .B1(new_n805), .B2(new_n807), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n296), .A2(new_n352), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n824), .A2(new_n666), .ZN(new_n988));
  OR4_X1    g802(.A1(new_n987), .A2(new_n988), .A3(new_n723), .A4(new_n771), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n985), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n981), .B1(new_n990), .B2(G953), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT127), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n981), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n793), .A2(new_n987), .A3(new_n834), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n983), .B(new_n780), .C1(new_n774), .C2(new_n775), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n986), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n330), .A2(G900), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n995), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n991), .A2(new_n994), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n994), .B1(new_n991), .B2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(G72));
  INV_X1    g818(.A(new_n713), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n990), .A2(new_n974), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n262), .A2(new_n245), .A3(new_n264), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n986), .A2(new_n974), .A3(new_n998), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n1008), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n1005), .A2(new_n865), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1013));
  NOR4_X1   g827(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .A4(new_n928), .ZN(G57));
endmodule


