//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  OR3_X1    g003(.A1(new_n189), .A2(KEYINPUT73), .A3(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n193));
  INV_X1    g007(.A(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(G146), .A3(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G128), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n203), .A2(KEYINPUT23), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(KEYINPUT23), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(new_n205), .C1(G119), .C2(new_n206), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n202), .A2(KEYINPUT71), .A3(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT71), .B1(new_n202), .B2(G128), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n208), .A2(new_n209), .B1(new_n202), .B2(G128), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT24), .B(G110), .Z(new_n211));
  AOI22_X1  g025(.A1(new_n207), .A2(G110), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n200), .A2(new_n212), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n207), .A2(G110), .B1(new_n210), .B2(new_n211), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n187), .A2(new_n197), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n199), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT22), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(G137), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n217), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT74), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(KEYINPUT25), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(KEYINPUT25), .ZN(new_n227));
  OR3_X1    g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G234), .ZN(new_n229));
  OAI21_X1  g043(.A(G217), .B1(new_n229), .B2(G902), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n224), .B2(new_n226), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(G902), .B1(new_n229), .B2(G217), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n234), .B(KEYINPUT75), .Z(new_n235));
  NOR2_X1   g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(G101), .ZN(new_n239));
  INV_X1    g053(.A(G237), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n218), .A3(G210), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n239), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT2), .B(G113), .Z(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n197), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n197), .A2(KEYINPUT64), .A3(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n253), .A2(new_n254), .A3(G128), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n249), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(G143), .B2(new_n197), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n206), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  INV_X1    g078(.A(G137), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT11), .A3(G134), .ZN(new_n266));
  INV_X1    g080(.A(G131), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(G137), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n264), .A2(new_n266), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n269), .A2(new_n270), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n263), .A2(G137), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n275), .B2(new_n268), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n261), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n264), .A2(new_n268), .A3(new_n266), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(KEYINPUT66), .B(new_n280), .C1(new_n271), .C2(new_n272), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n251), .A2(new_n252), .B1(new_n255), .B2(G146), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT0), .A3(G128), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n256), .A2(new_n249), .B1(KEYINPUT0), .B2(G128), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(KEYINPUT0), .B2(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT67), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n293), .B(new_n290), .C1(new_n283), .C2(new_n284), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n248), .B(new_n278), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n281), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n278), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n247), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n244), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n290), .B1(new_n283), .B2(new_n284), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n301), .A2(new_n247), .A3(new_n277), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n302), .B2(KEYINPUT28), .ZN(new_n303));
  INV_X1    g117(.A(new_n284), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n265), .A2(KEYINPUT11), .A3(G134), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT11), .B1(new_n265), .B2(G134), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(KEYINPUT65), .A3(new_n267), .A4(new_n268), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n269), .A2(new_n270), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT66), .B1(new_n310), .B2(new_n280), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n291), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n278), .A3(new_n248), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT69), .A3(new_n244), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n303), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n243), .B1(new_n299), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n295), .A2(new_n242), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n278), .A2(new_n318), .A3(new_n296), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n293), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n301), .A2(KEYINPUT67), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n277), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n322), .B2(new_n318), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n317), .B1(new_n323), .B2(new_n247), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n247), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n243), .B1(new_n322), .B2(new_n248), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n325), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n319), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n278), .B1(new_n292), .B2(new_n294), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(KEYINPUT30), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n329), .B(new_n325), .C1(new_n333), .C2(new_n248), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n330), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n302), .A2(new_n300), .A3(KEYINPUT28), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT69), .B1(new_n313), .B2(new_n244), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n295), .A2(new_n298), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(new_n244), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n329), .B1(new_n333), .B2(new_n248), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n345), .A2(new_n243), .B1(new_n346), .B2(KEYINPUT31), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n338), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n332), .A2(new_n247), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n295), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n315), .B1(new_n353), .B2(KEYINPUT28), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n243), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n242), .B1(new_n299), .B2(new_n315), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n295), .B(new_n243), .C1(new_n333), .C2(new_n248), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT70), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n299), .A2(new_n315), .A3(new_n243), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n355), .B1(new_n361), .B2(KEYINPUT70), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n357), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G472), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n237), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(KEYINPUT78), .A2(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT78), .A2(G107), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(G104), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G104), .A2(G107), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT3), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT3), .A3(G104), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OR4_X1    g191(.A1(KEYINPUT4), .A2(new_n373), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n374), .B1(new_n373), .B2(new_n377), .ZN(new_n379));
  AND2_X1   g193(.A1(KEYINPUT78), .A2(G107), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT78), .A2(G107), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n371), .B1(new_n382), .B2(G104), .ZN(new_n383));
  OAI211_X1 g197(.A(G101), .B(new_n376), .C1(new_n383), .C2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n384), .A3(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n385), .A3(new_n247), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n375), .A2(G104), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n374), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n376), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n374), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n202), .A2(G116), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(KEYINPUT5), .B2(new_n246), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n397), .A2(G113), .B1(new_n246), .B2(new_n245), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(G110), .B(G122), .Z(new_n401));
  OR2_X1    g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n401), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n261), .A2(new_n189), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n189), .B2(new_n291), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n218), .A2(G224), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT87), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n406), .B(new_n408), .Z(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n410), .A3(new_n401), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n394), .A2(new_n398), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT88), .A3(new_n399), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n401), .B(KEYINPUT8), .Z(new_n419));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n394), .A2(new_n420), .A3(new_n398), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n406), .A2(new_n413), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n416), .A2(new_n422), .A3(new_n423), .A4(new_n402), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n412), .A2(new_n424), .A3(new_n223), .ZN(new_n425));
  OAI21_X1  g239(.A(G210), .B1(G237), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT90), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n429), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n367), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G478), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(KEYINPUT15), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G116), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G122), .ZN(new_n437));
  INV_X1    g251(.A(G122), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G116), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n440), .A2(new_n382), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT96), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(KEYINPUT14), .A3(G122), .ZN(new_n443));
  OAI211_X1 g257(.A(G107), .B(new_n443), .C1(new_n440), .C2(KEYINPUT14), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT93), .B1(new_n206), .B2(G143), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n255), .A3(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n206), .A2(G143), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n448), .A2(new_n263), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n263), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n444), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT97), .B1(new_n442), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT96), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n441), .B(new_n454), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n450), .A2(new_n451), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .A4(new_n444), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT13), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n448), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n448), .A2(new_n461), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT94), .A4(KEYINPUT13), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n462), .A2(new_n449), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n440), .A2(new_n382), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n465), .A2(G134), .B1(new_n441), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n450), .B(KEYINPUT95), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT9), .B(G234), .Z(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(G217), .A3(new_n218), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n459), .B2(new_n469), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n223), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT98), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT98), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n223), .C1(new_n473), .C2(new_n475), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n435), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n434), .B1(new_n476), .B2(KEYINPUT98), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT99), .ZN(new_n483));
  INV_X1    g297(.A(G952), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G953), .ZN(new_n485));
  NAND2_X1  g299(.A1(G234), .A2(G237), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT21), .B(G898), .Z(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(G902), .A3(G953), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n240), .A2(new_n218), .A3(G214), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n255), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT17), .A3(G131), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(G131), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n494), .B(G143), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n267), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n198), .A2(new_n199), .A3(new_n496), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT18), .A2(G131), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n495), .B(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n215), .B1(new_n191), .B2(new_n197), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n390), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(new_n509), .A3(new_n506), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT92), .B(G475), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n497), .A2(new_n499), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n187), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n197), .B(new_n519), .C1(new_n191), .C2(new_n518), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n199), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n506), .A2(new_n521), .A3(KEYINPUT91), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT91), .B1(new_n506), .B2(new_n521), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n522), .A2(new_n523), .A3(new_n509), .ZN(new_n524));
  INV_X1    g338(.A(new_n512), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n516), .B(new_n223), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT20), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n523), .A2(new_n509), .ZN(new_n528));
  INV_X1    g342(.A(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n512), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n516), .A4(new_n223), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n493), .B(new_n515), .C1(new_n527), .C2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n482), .A2(new_n483), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n483), .B1(new_n482), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n432), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n471), .ZN(new_n538));
  OAI21_X1  g352(.A(G221), .B1(new_n538), .B2(G902), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT76), .Z(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G469), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n223), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n218), .A2(G227), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n194), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT77), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n546), .B(G110), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n285), .ZN(new_n549));
  INV_X1    g363(.A(new_n392), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n379), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n551), .A2(new_n261), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT83), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n257), .A2(KEYINPUT81), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n253), .A2(new_n256), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n259), .A2(KEYINPUT82), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT82), .ZN(new_n559));
  OAI21_X1  g373(.A(G128), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n286), .A2(new_n562), .A3(new_n254), .A4(G128), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n555), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n554), .B1(new_n564), .B2(new_n551), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n561), .A3(new_n563), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n394), .A2(new_n566), .A3(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n553), .B1(new_n568), .B2(new_n552), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n378), .A2(new_n385), .A3(new_n291), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT79), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n378), .A2(new_n385), .A3(new_n572), .A4(new_n291), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n549), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n394), .A2(new_n566), .A3(KEYINPUT83), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT83), .B1(new_n394), .B2(new_n566), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n552), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n553), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n549), .A2(new_n574), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n548), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n574), .A2(new_n578), .A3(new_n549), .A4(new_n579), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n551), .A2(new_n261), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n584), .A2(new_n281), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT12), .B1(new_n584), .B2(new_n285), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n582), .B(new_n547), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n543), .B1(new_n589), .B2(new_n542), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT85), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n582), .C1(new_n586), .C2(new_n587), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n548), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT86), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n580), .B2(new_n548), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n582), .A2(KEYINPUT86), .A3(new_n547), .ZN(new_n598));
  INV_X1    g412(.A(new_n575), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(G469), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n541), .B1(new_n590), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n537), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n365), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  OAI21_X1  g420(.A(G472), .B1(new_n336), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n348), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n602), .A4(new_n236), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n340), .A2(new_n347), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n223), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n348), .B1(new_n613), .B2(G472), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n614), .A2(KEYINPUT100), .A3(new_n236), .A4(new_n602), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n425), .A2(new_n426), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n412), .A2(new_n424), .A3(new_n223), .A4(new_n427), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n366), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n493), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n473), .A2(new_n475), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n470), .A2(KEYINPUT101), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n473), .A2(new_n475), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(KEYINPUT33), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G478), .B1(new_n628), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n527), .A2(new_n533), .ZN(new_n630));
  INV_X1    g444(.A(new_n515), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n622), .A2(new_n433), .A3(new_n223), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n621), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n616), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n630), .B(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n482), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n631), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n621), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n616), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(new_n221), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT103), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n217), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n233), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n232), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n604), .A2(new_n614), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT37), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G110), .ZN(G12));
  AOI21_X1  g469(.A(new_n349), .B1(new_n612), .B2(new_n337), .ZN(new_n656));
  AOI211_X1 g470(.A(KEYINPUT32), .B(new_n338), .C1(new_n340), .C2(new_n347), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n364), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n541), .B(new_n619), .C1(new_n601), .C2(new_n590), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n492), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n487), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n658), .A2(new_n659), .A3(new_n652), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT104), .B(G128), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G30));
  XOR2_X1   g481(.A(new_n662), .B(KEYINPUT39), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n602), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  AOI21_X1  g485(.A(new_n243), .B1(new_n327), .B2(new_n295), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n223), .B1(new_n353), .B2(new_n242), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n656), .B2(new_n657), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n430), .A2(new_n431), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT38), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n632), .B1(new_n480), .B2(new_n481), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n652), .A2(new_n367), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n671), .A2(new_n675), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  NOR2_X1   g495(.A1(new_n634), .A2(new_n663), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n658), .A2(new_n659), .A3(new_n652), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  XNOR2_X1  g498(.A(new_n589), .B(new_n542), .ZN(new_n685));
  INV_X1    g499(.A(new_n539), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n658), .A2(new_n635), .A3(new_n236), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n658), .A2(new_n643), .A3(new_n236), .A4(new_n687), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  OR2_X1    g506(.A1(new_n535), .A2(new_n536), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n685), .A2(new_n686), .A3(new_n619), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n658), .A2(new_n693), .A3(new_n652), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT105), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND2_X1  g511(.A1(new_n346), .A2(KEYINPUT31), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n354), .B2(new_n242), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n698), .B(KEYINPUT106), .C1(new_n242), .C2(new_n354), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n340), .A3(new_n702), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n703), .A2(new_n337), .B1(new_n613), .B2(G472), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n685), .A2(new_n686), .A3(new_n678), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n236), .A4(new_n620), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND4_X1  g521(.A1(new_n704), .A2(new_n652), .A3(new_n682), .A4(new_n694), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NAND3_X1  g523(.A1(new_n430), .A2(new_n366), .A3(new_n431), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n634), .A2(new_n710), .A3(new_n663), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n686), .B1(new_n590), .B2(new_n601), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n365), .A2(KEYINPUT42), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n658), .A2(new_n236), .A3(new_n711), .A4(new_n712), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT42), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  AND4_X1   g532(.A1(new_n658), .A2(new_n236), .A3(new_n664), .A4(new_n712), .ZN(new_n719));
  INV_X1    g533(.A(new_n710), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  AND2_X1   g536(.A1(new_n595), .A2(new_n600), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT107), .B(G469), .C1(new_n723), .C2(KEYINPUT45), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n595), .A2(KEYINPUT45), .A3(new_n600), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n595), .B2(new_n600), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n542), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n543), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT46), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n589), .A2(new_n542), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n686), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n629), .A2(new_n633), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n632), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT43), .ZN(new_n739));
  INV_X1    g553(.A(new_n614), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n652), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n710), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n736), .A2(new_n669), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n735), .B2(new_n686), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n732), .A2(new_n734), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT47), .B(new_n539), .C1(new_n749), .C2(new_n731), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n711), .ZN(new_n752));
  OR3_X1    g566(.A1(new_n752), .A2(new_n658), .A3(new_n236), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT108), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  OR2_X1    g569(.A1(new_n685), .A2(KEYINPUT117), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n685), .A2(KEYINPUT117), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n541), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n748), .A2(new_n750), .A3(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n704), .A2(new_n236), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(new_n488), .A3(new_n739), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT116), .B1(new_n761), .B2(new_n720), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n488), .A3(new_n739), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n763), .A2(new_n764), .A3(new_n710), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n677), .A2(new_n366), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n687), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n685), .A2(new_n710), .A3(new_n686), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(KEYINPUT118), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(KEYINPUT118), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n487), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n515), .B1(new_n527), .B2(new_n533), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n675), .A2(new_n237), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n737), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n739), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n704), .A2(new_n652), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n767), .A2(new_n771), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n761), .A2(new_n694), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n759), .B2(new_n766), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n780), .A4(new_n771), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n787), .A2(new_n485), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(new_n365), .A3(new_n739), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT48), .Z(new_n793));
  NAND2_X1  g607(.A1(new_n775), .A2(new_n777), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n634), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n791), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n713), .A2(new_n716), .B1(new_n720), .B2(new_n719), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n704), .A2(new_n682), .A3(new_n712), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n658), .A2(new_n602), .A3(new_n482), .A4(new_n662), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n640), .A2(new_n631), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n652), .A3(new_n720), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT109), .B1(new_n482), .B2(new_n632), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n776), .B(new_n804), .C1(new_n480), .C2(new_n481), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n634), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n493), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n806), .A2(new_n432), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n611), .A2(new_n615), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n605), .A3(new_n653), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n688), .A2(new_n691), .A3(new_n695), .A4(new_n706), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n797), .A2(new_n802), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT110), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n665), .A2(new_n708), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n652), .A2(new_n663), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n678), .A2(new_n619), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n712), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n675), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n683), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n665), .A2(new_n708), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n820), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n665), .A2(new_n683), .A3(new_n708), .A4(new_n819), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n823), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n813), .A2(new_n814), .A3(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n802), .A2(new_n797), .A3(new_n810), .A4(new_n811), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n815), .A2(new_n820), .A3(KEYINPUT52), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT113), .B1(new_n836), .B2(new_n831), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n833), .A2(KEYINPUT53), .A3(new_n835), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n829), .A2(new_n830), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n821), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n836), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n812), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT115), .B1(new_n851), .B2(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n839), .A2(new_n853), .A3(new_n814), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n846), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n845), .B1(new_n855), .B2(new_n842), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n796), .B(new_n844), .C1(new_n843), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n484), .A2(new_n218), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n677), .A2(new_n632), .A3(new_n737), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n540), .B1(new_n685), .B2(KEYINPUT49), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(KEYINPUT49), .B2(new_n685), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n777), .A3(new_n862), .A4(new_n366), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(G75));
  INV_X1    g678(.A(new_n846), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n851), .A2(KEYINPUT115), .A3(KEYINPUT53), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n853), .B1(new_n839), .B2(new_n814), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(G210), .A3(G902), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT120), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n855), .A2(new_n223), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(G210), .ZN(new_n873));
  XNOR2_X1  g687(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n404), .A2(new_n411), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n409), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n878), .B2(KEYINPUT122), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n878), .A2(KEYINPUT122), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n870), .A2(new_n873), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n218), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n869), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n884), .B2(new_n877), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n881), .A2(new_n885), .ZN(G51));
  NAND2_X1  g700(.A1(new_n581), .A2(new_n588), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n730), .A2(KEYINPUT57), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n855), .A2(new_n842), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT54), .B(new_n846), .C1(new_n852), .C2(new_n854), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n730), .A2(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n855), .A2(new_n223), .A3(new_n729), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n882), .B1(new_n893), .B2(new_n894), .ZN(G54));
  NAND3_X1  g709(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n512), .A3(new_n530), .ZN(new_n897));
  INV_X1    g711(.A(new_n882), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .A4(new_n531), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G60));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT59), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n889), .B2(new_n890), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n898), .B1(new_n903), .B2(new_n628), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n856), .A2(new_n843), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n841), .A2(new_n845), .A3(new_n842), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n907), .B2(new_n628), .ZN(G63));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT60), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n868), .A2(new_n650), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n222), .B(KEYINPUT124), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n855), .B2(new_n910), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n868), .A2(KEYINPUT123), .A3(new_n650), .A4(new_n911), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n914), .A2(new_n898), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n916), .A2(new_n898), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(new_n914), .A3(KEYINPUT61), .A4(new_n917), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(G66));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n810), .A2(new_n811), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT125), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n218), .ZN(new_n927));
  INV_X1    g741(.A(G224), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n490), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n924), .B2(new_n929), .ZN(new_n931));
  INV_X1    g745(.A(G898), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n875), .B1(new_n932), .B2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  AND3_X1   g748(.A1(new_n824), .A2(new_n683), .A3(new_n827), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n680), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n670), .A2(new_n710), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n365), .A2(new_n806), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n745), .A3(new_n753), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n218), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n519), .B1(new_n191), .B2(new_n518), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n323), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(G227), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n945), .B2(new_n660), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT127), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n736), .A2(new_n365), .A3(new_n669), .A4(new_n817), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n797), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n753), .A2(new_n950), .A3(new_n745), .A4(new_n935), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n218), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n660), .A2(G953), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n944), .B(new_n948), .C1(new_n954), .C2(new_n943), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n956));
  INV_X1    g770(.A(new_n943), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n940), .B2(new_n218), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n947), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n955), .A2(new_n959), .ZN(G72));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n940), .B2(new_n926), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n672), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n951), .B2(new_n926), .ZN(new_n965));
  INV_X1    g779(.A(new_n359), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n962), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n841), .A2(new_n966), .A3(new_n672), .A4(new_n968), .ZN(new_n969));
  NOR4_X1   g783(.A1(new_n964), .A2(new_n967), .A3(new_n882), .A4(new_n969), .ZN(G57));
endmodule


