//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1311, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AND2_X1   g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G244), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n215), .A2(G77), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(new_n213), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G250), .B(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G264), .B(G270), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n228), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT66), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G68), .Z(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  XNOR2_X1  g0042(.A(KEYINPUT3), .B(G33), .ZN(new_n243));
  INV_X1    g0043(.A(G1698), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n243), .A2(G222), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n243), .A2(G223), .A3(G1698), .ZN(new_n246));
  OAI211_X1 g0046(.A(new_n245), .B(new_n246), .C1(new_n202), .C2(new_n243), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n212), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  OAI21_X1  g0053(.A(G274), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(new_n205), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n254), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n205), .A2(new_n259), .B1(new_n212), .B2(new_n248), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(G226), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G200), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n251), .A2(new_n264), .A3(G190), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n253), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n206), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT68), .B1(G20), .B2(G33), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(G33), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n279), .A2(new_n280), .B1(new_n206), .B2(new_n201), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n271), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n206), .A3(G1), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n271), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n205), .B2(G20), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(new_n286), .B2(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n268), .B1(new_n269), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n269), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT72), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(KEYINPUT10), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n290), .B(new_n293), .C1(KEYINPUT10), .C2(new_n295), .ZN(new_n298));
  INV_X1    g0098(.A(new_n289), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n265), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(G179), .B2(new_n265), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n276), .A2(new_n286), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n280), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n271), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n271), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n283), .A2(G1), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G20), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(KEYINPUT69), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT69), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n284), .B2(new_n271), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n205), .A2(G20), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n312), .A2(new_n314), .A3(G68), .A4(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT11), .B(new_n271), .C1(new_n304), .C2(new_n305), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n284), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT12), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n308), .A2(new_n316), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  INV_X1    g0122(.A(G226), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n244), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n230), .A2(G1698), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n328), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n333), .A3(new_n250), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n262), .B1(G238), .B2(new_n263), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n334), .B2(new_n335), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n322), .B(G169), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n335), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(G179), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n342), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n322), .B1(new_n345), .B2(G169), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n321), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(new_n342), .A3(G190), .ZN(new_n349));
  INV_X1    g0149(.A(new_n321), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n279), .B1(new_n205), .B2(G20), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n285), .B1(new_n284), .B2(new_n279), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n274), .A2(new_n275), .ZN(new_n357));
  XNOR2_X1  g0157(.A(G58), .B(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(G159), .B1(new_n358), .B2(G20), .ZN(new_n359));
  OR2_X1    g0159(.A1(KEYINPUT3), .A2(G33), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n206), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n361), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n318), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n359), .B1(new_n366), .B2(KEYINPUT75), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT75), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n368), .B(new_n318), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n356), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n358), .A2(G20), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n276), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n309), .B1(new_n374), .B2(KEYINPUT16), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n355), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n261), .A2(new_n256), .ZN(new_n377));
  INV_X1    g0177(.A(new_n254), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n249), .A2(G232), .A3(new_n255), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G223), .A2(G1698), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n323), .B2(G1698), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n243), .B1(G33), .B2(G87), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n379), .B(new_n381), .C1(new_n384), .C2(new_n249), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G169), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n323), .A2(G1698), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n387), .B1(G223), .B2(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n250), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n391), .A2(G179), .A3(new_n379), .A4(new_n381), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT18), .B1(new_n376), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n326), .A2(new_n327), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n396), .B2(new_n206), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n326), .A2(new_n327), .A3(new_n363), .A4(G20), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n373), .B1(new_n399), .B2(new_n368), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n366), .A2(KEYINPUT75), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n271), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n354), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n393), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n385), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n391), .A2(new_n410), .A3(new_n379), .A4(new_n381), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n354), .C1(new_n402), .C2(new_n404), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n376), .A2(KEYINPUT17), .A3(new_n412), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n395), .A2(new_n407), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT71), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n279), .B1(new_n274), .B2(new_n275), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n280), .B1(new_n206), .B2(new_n202), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n271), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n312), .A2(new_n314), .A3(G77), .A4(new_n315), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n284), .A2(new_n202), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(G232), .B(new_n244), .C1(new_n326), .C2(new_n327), .ZN(new_n426));
  OAI211_X1 g0226(.A(G238), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n427));
  INV_X1    g0227(.A(G107), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(new_n427), .C1(new_n428), .C2(new_n243), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n250), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n377), .A2(new_n378), .B1(new_n263), .B2(new_n215), .ZN(new_n431));
  AOI21_X1  g0231(.A(G169), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n418), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n431), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n300), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT71), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT70), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n434), .B2(G179), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT70), .A4(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n433), .A2(new_n437), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n436), .B1(G200), .B2(new_n434), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n410), .B2(new_n434), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR4_X1   g0245(.A1(new_n303), .A2(new_n352), .A3(new_n417), .A4(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(G244), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT78), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT78), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n243), .A2(new_n449), .A3(G244), .A4(G1698), .ZN(new_n450));
  OR2_X1    g0250(.A1(KEYINPUT79), .A2(G116), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT79), .A2(G116), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n273), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n243), .A2(G238), .A3(new_n244), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n448), .A2(new_n450), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n250), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n205), .A2(G45), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n249), .A2(G250), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n254), .B2(new_n458), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n440), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n457), .B2(new_n461), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT80), .B(new_n460), .C1(new_n456), .C2(new_n250), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n300), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT19), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n206), .B1(new_n329), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G87), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n428), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n243), .A2(new_n206), .A3(G68), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n470), .B1(new_n280), .B2(new_n473), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n271), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n420), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n311), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n205), .A2(G33), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n285), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n481), .B(new_n484), .C1(new_n420), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n466), .A2(new_n469), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n463), .A2(G190), .A3(new_n465), .ZN(new_n489));
  OAI21_X1  g0289(.A(G200), .B1(new_n467), .B2(new_n468), .ZN(new_n490));
  INV_X1    g0290(.A(new_n486), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n481), .A2(new_n484), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n451), .A2(G20), .A3(new_n452), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n206), .C1(G33), .C2(new_n473), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n271), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n312), .A2(new_n314), .A3(G116), .A4(new_n485), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n451), .A2(new_n452), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G20), .A3(new_n310), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n243), .A2(G264), .A3(G1698), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n396), .A2(G303), .ZN(new_n509));
  OAI211_X1 g0309(.A(G257), .B(new_n244), .C1(new_n326), .C2(new_n327), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT5), .B(G41), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n258), .A2(G1), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n512), .A2(new_n513), .B1(new_n212), .B2(new_n248), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n511), .A2(new_n250), .B1(G270), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n458), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n378), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n507), .A2(G179), .A3(new_n515), .A4(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n511), .A2(new_n250), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n514), .A2(G270), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n520), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n515), .A2(G190), .A3(new_n520), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n300), .B1(new_n515), .B2(new_n520), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT82), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(KEYINPUT21), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n529), .A2(new_n507), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n529), .B2(new_n507), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n521), .B(new_n528), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n514), .A2(G264), .B1(new_n378), .B2(new_n519), .ZN(new_n536));
  OAI211_X1 g0336(.A(G257), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n537));
  OAI211_X1 g0337(.A(G250), .B(new_n244), .C1(new_n326), .C2(new_n327), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G294), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n250), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(new_n541), .A3(G179), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n514), .A2(G264), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n520), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n541), .A2(KEYINPUT83), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n540), .A2(new_n546), .A3(new_n250), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n542), .B1(new_n548), .B2(new_n300), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n206), .B(G87), .C1(new_n326), .C2(new_n327), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT22), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n243), .A2(new_n552), .A3(new_n206), .A4(G87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n206), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n428), .A2(KEYINPUT23), .A3(G20), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n453), .A2(new_n206), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n555), .B1(new_n554), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n271), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n311), .B2(G107), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n428), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n491), .A2(G107), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n549), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n540), .A2(new_n546), .A3(new_n250), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n546), .B1(new_n540), .B2(new_n250), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n410), .B(new_n536), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n536), .A2(new_n541), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n408), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n562), .A3(new_n566), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(new_n244), .C1(new_n326), .C2(new_n327), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n243), .A2(KEYINPUT4), .A3(G244), .A4(new_n244), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(new_n579), .A3(new_n498), .ZN(new_n580));
  OAI211_X1 g0380(.A(G250), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n249), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT77), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n514), .B2(G257), .ZN(new_n585));
  AND2_X1   g0385(.A1(KEYINPUT5), .A2(G41), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n513), .B1(new_n586), .B2(new_n516), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G257), .A3(new_n249), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n520), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n300), .B1(new_n583), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT76), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n581), .B(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n578), .A2(new_n579), .A3(new_n498), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n250), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n514), .A2(new_n584), .A3(G257), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n378), .B2(new_n519), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n598), .A3(new_n440), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n600), .A2(new_n473), .A3(G107), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n206), .B1(new_n202), .B2(new_n276), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n428), .B1(new_n364), .B2(new_n365), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n271), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n284), .A2(new_n473), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n491), .A2(G97), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n591), .A2(new_n599), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(G200), .B1(new_n583), .B2(new_n590), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n607), .B1(new_n486), .B2(new_n473), .ZN(new_n612));
  INV_X1    g0412(.A(new_n605), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n602), .A2(new_n600), .ZN(new_n614));
  INV_X1    g0414(.A(new_n601), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(G20), .B1(G77), .B2(new_n357), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n618), .B2(new_n271), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n595), .A2(new_n598), .A3(G190), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n611), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n568), .A2(new_n575), .A3(new_n610), .A4(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n446), .A2(new_n496), .A3(new_n535), .A4(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n446), .ZN(new_n624));
  INV_X1    g0424(.A(new_n610), .ZN(new_n625));
  AND4_X1   g0425(.A1(KEYINPUT26), .A2(new_n488), .A3(new_n495), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n487), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n467), .A2(new_n468), .A3(G179), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n462), .A2(new_n300), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n466), .A2(KEYINPUT84), .A3(new_n631), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n481), .A2(new_n637), .A3(new_n484), .A4(new_n492), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n462), .A2(G200), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(new_n489), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n635), .A2(new_n610), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n627), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n630), .A2(new_n629), .A3(new_n632), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT84), .B1(new_n466), .B2(new_n631), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n487), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n515), .A2(G179), .A3(new_n520), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n522), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n525), .A2(G169), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n522), .A2(new_n649), .B1(new_n530), .B2(KEYINPUT21), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n529), .A2(new_n507), .A3(new_n531), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n549), .A2(new_n567), .A3(KEYINPUT86), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT86), .B1(new_n549), .B2(new_n567), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n639), .A2(new_n489), .A3(new_n640), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n575), .A2(new_n610), .A3(new_n621), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n646), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n646), .A2(KEYINPUT87), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT87), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n635), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n624), .B1(new_n643), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n395), .A2(new_n407), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n347), .A2(new_n442), .ZN(new_n666));
  INV_X1    g0466(.A(new_n351), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n413), .A2(new_n414), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT17), .B1(new_n376), .B2(new_n412), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n297), .A2(new_n298), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n302), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n663), .A2(new_n673), .ZN(G369));
  NOR3_X1   g0474(.A1(new_n283), .A2(G1), .A3(G20), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT27), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G213), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n675), .B2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT88), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n677), .A2(new_n679), .A3(new_n683), .A4(G343), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n652), .A2(new_n522), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n535), .B1(new_n522), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n692), .A3(G330), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n568), .A2(new_n575), .ZN(new_n695));
  INV_X1    g0495(.A(new_n567), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n686), .ZN(new_n697));
  INV_X1    g0497(.A(new_n568), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n685), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n652), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n695), .A2(new_n702), .A3(new_n686), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n653), .A2(new_n654), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n685), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n701), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n209), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n474), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n214), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n463), .A2(new_n465), .ZN(new_n715));
  INV_X1    g0515(.A(new_n542), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n515), .A3(new_n595), .A4(new_n598), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n595), .A2(new_n598), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n515), .A2(G179), .A3(new_n536), .A4(new_n541), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n463), .A4(new_n465), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n536), .B2(new_n541), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n719), .A2(new_n462), .A3(new_n525), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n685), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n496), .A2(new_n622), .A3(new_n535), .A4(new_n686), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n652), .A2(new_n568), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n646), .A2(new_n656), .A3(new_n657), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT26), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n496), .A2(new_n736), .A3(new_n625), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n735), .A2(new_n659), .A3(new_n661), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n642), .A2(new_n736), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT29), .B(new_n686), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n635), .B(KEYINPUT87), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n646), .A2(new_n625), .A3(new_n656), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT26), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n742), .A2(new_n744), .A3(new_n735), .A4(new_n737), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT90), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT29), .A4(new_n686), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n626), .B1(new_n743), .B2(new_n736), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n686), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n733), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n713), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(new_n694), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n283), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n205), .B1(new_n757), .B2(G45), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n709), .A2(KEYINPUT91), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT91), .ZN(new_n760));
  INV_X1    g0560(.A(new_n758), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n708), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n756), .B(new_n763), .C1(G330), .C2(new_n689), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n253), .B1(G20), .B2(new_n300), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n440), .A2(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n206), .A2(G190), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT96), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT96), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G58), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n206), .A2(new_n410), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n767), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n771), .A2(new_n202), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G159), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n408), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n243), .B1(new_n783), .B2(new_n472), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n768), .A2(new_n782), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(G107), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n410), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n780), .A2(KEYINPUT32), .B1(new_n789), .B2(G50), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n206), .B1(new_n777), .B2(G190), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n473), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n788), .A2(G190), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(G68), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n781), .A2(new_n787), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n776), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n779), .A2(G329), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n783), .C1(new_n799), .C2(new_n774), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n771), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  INV_X1    g0603(.A(new_n793), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT33), .B(G317), .Z(new_n805));
  OAI221_X1 g0605(.A(new_n396), .B1(new_n785), .B2(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n789), .A2(G326), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n791), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n800), .A2(new_n802), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n766), .B1(new_n796), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n707), .A2(new_n243), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G45), .B2(new_n214), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(KEYINPUT95), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(KEYINPUT95), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n258), .C2(new_n241), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT93), .ZN(new_n817));
  NAND2_X1  g0617(.A1(G355), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(G355), .A2(new_n817), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n209), .A2(new_n243), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(G116), .B2(new_n209), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT94), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n816), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n766), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n763), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n828), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n811), .B(new_n830), .C1(new_n689), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n765), .A2(new_n832), .A3(new_n833), .ZN(G396));
  INV_X1    g0634(.A(new_n774), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(G143), .B1(G137), .B2(new_n789), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n277), .B2(new_n804), .C1(new_n372), .C2(new_n771), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  INV_X1    g0638(.A(new_n783), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n396), .B1(new_n839), .B2(G50), .ZN(new_n840));
  INV_X1    g0640(.A(new_n791), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G58), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n786), .A2(G68), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n779), .A2(G132), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n789), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n798), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n792), .B(new_n847), .C1(G283), .C2(new_n793), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n785), .A2(new_n472), .B1(new_n778), .B2(new_n801), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G294), .B2(new_n835), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(new_n505), .C2(new_n771), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n396), .B1(new_n783), .B2(new_n428), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT98), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n838), .A2(new_n845), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n766), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n766), .A2(new_n826), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n763), .B1(new_n202), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n685), .A2(new_n436), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n685), .B2(new_n436), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n442), .A2(new_n861), .A3(new_n444), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n442), .B2(new_n444), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n855), .B(new_n857), .C1(new_n865), .C2(new_n827), .ZN(new_n866));
  INV_X1    g0666(.A(new_n763), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n864), .A2(new_n685), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n662), .B2(new_n643), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n751), .B2(new_n864), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n867), .B1(new_n872), .B2(new_n732), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n732), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n866), .B1(new_n874), .B2(new_n875), .ZN(G384));
  INV_X1    g0676(.A(G116), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n877), .B(new_n213), .C1(new_n616), .C2(KEYINPUT35), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT35), .B2(new_n616), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT36), .ZN(new_n880));
  OAI21_X1  g0680(.A(G77), .B1(new_n772), .B2(new_n318), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n881), .A2(new_n214), .B1(G50), .B2(new_n318), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(G1), .A3(new_n283), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT100), .Z(new_n885));
  OAI21_X1  g0685(.A(new_n413), .B1(new_n376), .B2(new_n394), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n376), .A2(new_n680), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n405), .A2(new_n393), .ZN(new_n889));
  INV_X1    g0689(.A(new_n680), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n405), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n892), .A4(new_n413), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n417), .A2(new_n887), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT39), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n356), .B1(new_n366), .B2(new_n373), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n403), .A3(new_n271), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n900), .A2(new_n901), .A3(new_n354), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n900), .B2(new_n354), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n386), .A2(new_n392), .A3(new_n680), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n413), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n893), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n902), .A2(new_n903), .A3(new_n680), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n417), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT102), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n893), .A2(new_n907), .B1(new_n417), .B2(new_n909), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n898), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT39), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(G169), .B1(new_n337), .B2(new_n338), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT14), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n343), .A3(new_n339), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n321), .A3(new_n686), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n893), .ZN(new_n927));
  INV_X1    g0727(.A(new_n903), .ZN(new_n928));
  INV_X1    g0728(.A(new_n904), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n900), .A2(new_n901), .A3(new_n354), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n892), .B1(new_n931), .B2(new_n413), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n909), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n668), .A2(new_n669), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n664), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n897), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n911), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n321), .A2(new_n685), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n347), .A2(new_n351), .A3(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n321), .B(new_n685), .C1(new_n923), .C2(new_n667), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n442), .A2(new_n685), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n938), .B(new_n942), .C1(new_n870), .C2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n664), .A2(new_n890), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n926), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n945), .B1(new_n920), .B2(new_n925), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(KEYINPUT103), .A3(new_n944), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n624), .B1(new_n751), .B2(new_n752), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n673), .B1(new_n748), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n896), .A2(new_n897), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n913), .A2(new_n915), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n864), .B1(new_n940), .B2(new_n941), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n731), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT104), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n731), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n957), .A2(new_n960), .A3(KEYINPUT40), .A4(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n731), .B(new_n958), .C1(new_n917), .C2(new_n918), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT40), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n446), .A2(new_n731), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(G330), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n955), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n205), .B2(new_n757), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n955), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n885), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT105), .Z(G367));
  OAI211_X1 g0776(.A(new_n697), .B(new_n699), .C1(new_n652), .C2(new_n685), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n977), .A2(new_n703), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n691), .A2(new_n978), .A3(new_n693), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n703), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n692), .B1(new_n689), .B2(G330), .ZN(new_n981));
  INV_X1    g0781(.A(G330), .ZN(new_n982));
  AOI211_X1 g0782(.A(KEYINPUT89), .B(new_n982), .C1(new_n687), .C2(new_n688), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n754), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT112), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n754), .A2(KEYINPUT112), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n701), .A2(KEYINPUT111), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n610), .A2(new_n621), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n609), .A2(new_n685), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n992), .A2(new_n993), .B1(new_n625), .B2(new_n685), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n705), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT44), .Z(new_n996));
  NOR2_X1   g0796(.A1(new_n705), .A2(new_n994), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n991), .B(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n989), .A2(new_n990), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n754), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n708), .B(KEYINPUT41), .Z(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n761), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n635), .A2(new_n641), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n636), .A2(new_n638), .A3(new_n685), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n742), .B2(new_n1007), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT106), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT106), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n703), .A2(new_n994), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT42), .Z(new_n1015));
  NAND3_X1  g0815(.A1(new_n992), .A2(new_n698), .A3(new_n993), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1016), .A2(KEYINPUT108), .A3(new_n610), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT108), .B1(new_n1016), .B2(new_n610), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1017), .A2(new_n1018), .A3(new_n685), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1012), .A2(new_n1013), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT109), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1020), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1010), .A2(KEYINPUT43), .A3(new_n1011), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT110), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n1024), .A2(KEYINPUT110), .A3(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n701), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1029), .A2(new_n994), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1026), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1024), .A2(KEYINPUT110), .A3(new_n1025), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n1030), .A3(new_n1023), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n831), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n812), .A2(new_n227), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n829), .C1(new_n209), .C2(new_n420), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n771), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(G50), .ZN(new_n1042));
  INV_X1    g0842(.A(G137), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n785), .A2(new_n202), .B1(new_n778), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G58), .B2(new_n839), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n243), .B1(new_n774), .B2(new_n277), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G159), .B2(new_n793), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n791), .A2(new_n318), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n789), .B2(G143), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1042), .A2(new_n1045), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n839), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n428), .B2(new_n791), .C1(new_n798), .C2(new_n774), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G283), .B2(new_n1041), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT46), .B1(new_n839), .B2(new_n504), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G294), .B2(new_n793), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(new_n801), .C2(new_n846), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n785), .A2(new_n473), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n243), .B(new_n1057), .C1(G317), .C2(new_n779), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT113), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n1050), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT47), .Z(new_n1061));
  INV_X1    g0861(.A(new_n766), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n867), .B(new_n1040), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1005), .A2(new_n1037), .B1(new_n1038), .B2(new_n1063), .ZN(G387));
  NAND3_X1  g0864(.A1(new_n697), .A2(new_n699), .A3(new_n828), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n710), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n209), .A3(new_n243), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(G107), .B2(new_n209), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n707), .B(new_n243), .C1(new_n233), .C2(G45), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n258), .B1(new_n318), .B2(new_n202), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1066), .B2(KEYINPUT114), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n279), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1072), .A2(KEYINPUT50), .A3(new_n286), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT50), .B1(new_n1072), .B2(new_n286), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1071), .B1(KEYINPUT114), .B2(new_n1066), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1068), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n829), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n867), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n396), .B(new_n1057), .C1(G159), .C2(new_n789), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n791), .A2(new_n420), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n793), .B2(new_n1072), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1041), .A2(G68), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n783), .A2(new_n202), .B1(new_n778), .B2(new_n277), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G50), .B2(new_n835), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n243), .B1(new_n779), .B2(G326), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n783), .A2(new_n808), .B1(new_n791), .B2(new_n803), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n835), .A2(G317), .B1(G311), .B2(new_n793), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n799), .B2(new_n846), .C1(new_n798), .C2(new_n771), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT49), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1086), .B1(new_n505), .B2(new_n785), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1085), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1078), .B1(new_n1096), .B2(new_n766), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n986), .A2(new_n761), .B1(new_n1065), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n708), .B1(new_n754), .B2(new_n986), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT112), .B1(new_n754), .B2(new_n986), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n741), .A2(new_n747), .B1(new_n752), .B2(new_n751), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1101), .A2(new_n985), .A3(new_n988), .A4(new_n733), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1098), .B1(new_n1099), .B2(new_n1103), .ZN(G393));
  XNOR2_X1  g0904(.A(new_n999), .B(new_n701), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1001), .A2(new_n1106), .A3(new_n708), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT116), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1001), .A2(new_n1106), .A3(new_n1109), .A4(new_n708), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n835), .A2(G311), .B1(G317), .B2(new_n789), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT52), .Z(new_n1113));
  OAI22_X1  g0913(.A1(new_n783), .A2(new_n803), .B1(new_n778), .B2(new_n799), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n243), .B(new_n1114), .C1(G107), .C2(new_n786), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1041), .A2(G294), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n841), .A2(new_n504), .B1(G303), .B2(new_n793), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n846), .A2(new_n277), .B1(new_n774), .B2(new_n372), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n783), .A2(new_n318), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n243), .B1(new_n785), .B2(new_n472), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G143), .C2(new_n779), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1041), .A2(new_n1072), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n791), .A2(new_n202), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n793), .B2(G50), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1062), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n812), .A2(new_n237), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1077), .B1(G97), .B2(new_n707), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n763), .B(new_n1128), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT115), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n994), .A2(new_n828), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1105), .B2(new_n758), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1111), .A2(new_n1136), .ZN(G390));
  NAND3_X1  g0937(.A1(new_n733), .A2(new_n865), .A3(new_n942), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n942), .B1(new_n870), .B2(new_n943), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n920), .B1(new_n1140), .B2(new_n924), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n957), .A2(new_n924), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n686), .B(new_n865), .C1(new_n738), .C2(new_n739), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n943), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1145), .B2(new_n942), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n942), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1142), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT39), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n937), .B2(new_n911), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT102), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n1153));
  AND4_X1   g0953(.A1(KEYINPUT102), .A2(new_n908), .A3(KEYINPUT38), .A4(new_n910), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1155), .B2(new_n898), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n942), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n868), .B1(new_n749), .B2(new_n750), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n1144), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1156), .B1(new_n1159), .B2(new_n925), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1150), .A2(new_n1160), .A3(new_n1138), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1147), .A2(new_n761), .A3(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT117), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n624), .A2(new_n732), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n673), .B(new_n1164), .C1(new_n748), .C2(new_n953), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1157), .B1(new_n732), .B2(new_n864), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1138), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1158), .A2(new_n1144), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1138), .A2(new_n1144), .A3(new_n1166), .A4(new_n1143), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1138), .B1(new_n1150), .B2(new_n1160), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1141), .A2(new_n1146), .A3(new_n1139), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1147), .A2(new_n1165), .A3(new_n1161), .A4(new_n1171), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n708), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n843), .B1(new_n808), .B2(new_n778), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G116), .B2(new_n835), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n243), .B(new_n1125), .C1(G87), .C2(new_n839), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G107), .A2(new_n793), .B1(new_n789), .B2(G283), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1041), .A2(G97), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n783), .A2(new_n277), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT53), .ZN(new_n1185));
  INV_X1    g0985(.A(G128), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1184), .A2(new_n1185), .B1(new_n1186), .B2(new_n846), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1185), .B2(new_n1184), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n778), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n243), .B1(new_n785), .B2(new_n286), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G132), .C2(new_n835), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT54), .B(G143), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1041), .A2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n841), .A2(G159), .B1(G137), .B2(new_n793), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1188), .A2(new_n1192), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1062), .B1(new_n1183), .B2(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n763), .B(new_n1198), .C1(new_n279), .C2(new_n856), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n920), .B2(new_n827), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1163), .A2(new_n1177), .A3(new_n1200), .ZN(G378));
  INV_X1    g1001(.A(KEYINPUT120), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1164), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n954), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1174), .A2(new_n1173), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n1171), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n982), .B1(new_n964), .B2(new_n965), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n299), .A2(new_n680), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT55), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n303), .A2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1211));
  INV_X1    g1011(.A(new_n1209), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n297), .A2(new_n298), .A3(new_n302), .A4(new_n1212), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n963), .A2(new_n1207), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n963), .B2(new_n1207), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n950), .A2(KEYINPUT103), .A3(new_n944), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT103), .B1(new_n950), .B2(new_n944), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n963), .A2(new_n1207), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1216), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n963), .A2(new_n1207), .A3(new_n1216), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n949), .A3(new_n951), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1222), .A2(new_n1228), .A3(KEYINPUT57), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1202), .B1(new_n1206), .B2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1222), .A2(new_n1228), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1176), .A2(new_n1165), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1231), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT119), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n949), .A2(new_n1235), .A3(new_n951), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1227), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1219), .A2(new_n949), .A3(new_n1235), .A4(new_n951), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1237), .A2(new_n1238), .B1(new_n1176), .B2(new_n1165), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n708), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1234), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1216), .A2(new_n826), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n785), .A2(new_n772), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n774), .A2(new_n428), .B1(new_n778), .B2(new_n803), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n1041), .C2(new_n482), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n396), .A2(new_n257), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1246), .B(new_n1048), .C1(G77), .C2(new_n839), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G97), .A2(new_n793), .B1(new_n789), .B2(G116), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT58), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G50), .B1(new_n273), .B2(new_n257), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1249), .A2(new_n1250), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n846), .A2(new_n1189), .B1(new_n791), .B2(new_n277), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n793), .A2(G132), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n774), .B2(new_n1186), .C1(new_n783), .C2(new_n1193), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1253), .B(new_n1255), .C1(G137), .C2(new_n1041), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT59), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n273), .B(new_n257), .C1(new_n785), .C2(new_n372), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G124), .B2(new_n779), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1252), .B1(new_n1250), .B2(new_n1249), .C1(new_n1258), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n766), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n856), .A2(new_n286), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1242), .A2(new_n867), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n761), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1241), .A2(new_n1268), .ZN(G375));
  AND2_X1   g1069(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1204), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1172), .A3(new_n1004), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT121), .Z(new_n1273));
  NAND2_X1  g1073(.A1(new_n1157), .A2(new_n826), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT122), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n504), .A2(new_n793), .B1(new_n789), .B2(G294), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n771), .B2(new_n428), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT123), .Z(new_n1278));
  AOI22_X1  g1078(.A1(G97), .A2(new_n839), .B1(new_n835), .B2(G283), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n798), .B2(new_n778), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n396), .B1(new_n785), .B2(new_n202), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(new_n1278), .A2(new_n1080), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n396), .B(new_n1243), .C1(G132), .C2(new_n789), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1041), .A2(G150), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(G50), .A2(new_n841), .B1(new_n1194), .B2(new_n793), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n783), .A2(new_n372), .B1(new_n778), .B2(new_n1186), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(G137), .B2(new_n835), .ZN(new_n1287));
  AND4_X1   g1087(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n766), .B1(new_n1282), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n763), .B1(new_n318), .B2(new_n856), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1275), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1171), .B2(new_n761), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1273), .A2(new_n1292), .ZN(new_n1293));
  XOR2_X1   g1093(.A(new_n1293), .B(KEYINPUT124), .Z(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(G381));
  INV_X1    g1095(.A(G375), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1135), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1297));
  INV_X1    g1097(.A(G384), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1038), .A2(new_n1063), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1030), .B1(new_n1035), .B2(new_n1023), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n754), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1103), .B2(new_n1000), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n758), .B1(new_n1304), .B2(new_n1003), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1299), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G378), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(G393), .A2(G396), .ZN(new_n1308));
  AND4_X1   g1108(.A1(new_n1298), .A2(new_n1306), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .A4(new_n1309), .ZN(G407));
  NAND3_X1  g1110(.A1(new_n1296), .A2(new_n681), .A3(new_n1307), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(G407), .A2(G213), .A3(new_n1311), .ZN(G409));
  OAI211_X1 g1112(.A(G378), .B(new_n1268), .C1(new_n1234), .C2(new_n1240), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1222), .A2(new_n1228), .A3(new_n761), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1265), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1239), .A2(new_n1004), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(KEYINPUT125), .A3(new_n1265), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1307), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1313), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n678), .A2(G343), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT60), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1271), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n708), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1271), .B2(new_n1172), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1292), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1298), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1292), .B(G384), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1323), .A2(G2897), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1333), .B(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(G393), .A2(G396), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1337), .A2(new_n1308), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1306), .A2(G390), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(G387), .A2(new_n1297), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT126), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1339), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  AOI211_X1 g1144(.A(KEYINPUT126), .B(new_n1338), .C1(new_n1340), .C2(new_n1341), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1333), .ZN(new_n1347));
  AND4_X1   g1147(.A1(KEYINPUT63), .A2(new_n1322), .A3(new_n1324), .A4(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1323), .B1(new_n1313), .B2(new_n1321), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT63), .B1(new_n1349), .B2(new_n1347), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1306), .A2(G390), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(G387), .A2(new_n1297), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1343), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1338), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1342), .A2(new_n1343), .A3(new_n1339), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1336), .B(new_n1346), .C1(new_n1351), .C2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT127), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1325), .A2(new_n1335), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT61), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1359), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1322), .A2(new_n1324), .A3(new_n1347), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(KEYINPUT62), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1349), .A2(new_n1365), .A3(new_n1347), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1357), .B1(new_n1362), .B2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1358), .A2(new_n1368), .ZN(G405));
  NAND2_X1  g1169(.A1(G375), .A2(new_n1307), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1370), .A2(new_n1313), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(new_n1347), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1370), .A2(new_n1313), .A3(new_n1333), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(new_n1357), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1372), .A2(new_n1355), .A3(new_n1356), .A4(new_n1373), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1375), .A2(new_n1376), .ZN(G402));
endmodule


