//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n232), .A2(G50), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n235), .A2(new_n207), .ZN(new_n236));
  AND2_X1   g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR4_X1   g0037(.A1(new_n213), .A2(new_n229), .A3(new_n230), .A4(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  INV_X1    g0052(.A(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT67), .B(G50), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n251), .B(new_n256), .ZN(G351));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n207), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n221), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n235), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n261), .A2(KEYINPUT77), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT11), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT73), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n272), .B2(new_n263), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n206), .A2(G20), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n235), .A4(new_n262), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n273), .A2(G68), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT78), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT11), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n266), .A2(new_n278), .A3(new_n267), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(new_n215), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT12), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n269), .A2(new_n277), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G274), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(new_n216), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(G232), .A4(G1698), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G97), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT75), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n296), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G226), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT3), .B(G33), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n305), .A2(KEYINPUT75), .A3(G226), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n292), .B(new_n293), .C1(new_n307), .C2(new_n285), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n306), .ZN(new_n309));
  INV_X1    g0109(.A(new_n299), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n285), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT13), .B1(new_n311), .B2(new_n291), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n312), .A2(G190), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n282), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT76), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n308), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT76), .B(KEYINPUT13), .C1(new_n311), .C2(new_n291), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G200), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(G169), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT14), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n316), .A2(new_n323), .A3(G169), .A4(new_n317), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n312), .A2(new_n308), .A3(G179), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n320), .B1(new_n282), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n263), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT8), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n329), .A2(new_n330), .A3(G58), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n260), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n272), .A2(new_n202), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n328), .A2(new_n274), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n202), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  INV_X1    g0142(.A(new_n288), .ZN(new_n343));
  INV_X1    g0143(.A(new_n290), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(G226), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n285), .B1(new_n301), .B2(new_n221), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G222), .A2(G1698), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT69), .B(G223), .Z(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(G1698), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(new_n301), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n341), .B1(new_n342), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(KEYINPUT71), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n345), .A2(new_n355), .A3(new_n350), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n341), .B(KEYINPUT9), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(G200), .B2(new_n351), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n359), .A2(new_n362), .A3(KEYINPUT74), .A4(KEYINPUT10), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n364));
  OR2_X1    g0164(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n365));
  INV_X1    g0165(.A(new_n362), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n358), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n288), .B1(new_n290), .B2(new_n222), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n305), .A2(G232), .A3(new_n302), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n305), .A2(G238), .A3(G1698), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n371), .C1(new_n223), .C2(new_n305), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n355), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G169), .B2(new_n374), .ZN(new_n376));
  INV_X1    g0176(.A(new_n258), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n332), .A2(new_n377), .B1(new_n207), .B2(new_n221), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(KEYINPUT72), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT15), .B(G87), .Z(new_n380));
  AOI22_X1  g0180(.A1(new_n378), .A2(KEYINPUT72), .B1(new_n334), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n328), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n273), .A2(G77), .A3(new_n274), .A4(new_n275), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G77), .B2(new_n271), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n374), .A2(G190), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n385), .B(new_n388), .C1(new_n389), .C2(new_n374), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n327), .A2(new_n357), .A3(new_n368), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n305), .B2(G20), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n294), .A2(G33), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT7), .B(new_n207), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n215), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n253), .A2(new_n215), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n258), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n393), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT79), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n283), .B2(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n294), .A2(KEYINPUT79), .A3(G33), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n296), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(new_n394), .A3(new_n207), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n394), .B1(new_n411), .B2(new_n207), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT16), .B(new_n407), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT81), .B(new_n393), .C1(new_n399), .C2(new_n403), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n406), .A2(new_n263), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n333), .A2(new_n339), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n333), .B2(new_n272), .ZN(new_n419));
  OR2_X1    g0219(.A1(G223), .A2(G1698), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(G226), .B2(new_n302), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n411), .A2(new_n421), .B1(new_n283), .B2(new_n217), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n373), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n288), .B1(new_n290), .B2(new_n240), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n425), .A3(new_n360), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n373), .B2(new_n422), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(G200), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n417), .A2(KEYINPUT84), .A3(new_n419), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT83), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n417), .A2(new_n433), .A3(new_n419), .A4(new_n428), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT82), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n427), .B2(new_n355), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G169), .B2(new_n427), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n427), .A2(new_n438), .A3(new_n355), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n417), .A2(new_n419), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n392), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n328), .B(new_n271), .C1(G1), .C2(new_n283), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n380), .ZN(new_n453));
  INV_X1    g0253(.A(new_n380), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n272), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n260), .A2(KEYINPUT19), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n217), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n298), .A2(new_n207), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n461), .B2(KEYINPUT19), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n409), .A2(new_n410), .A3(new_n296), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT86), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n207), .A4(G68), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n409), .A2(new_n410), .A3(new_n207), .A4(new_n296), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT86), .B1(new_n466), .B2(new_n215), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n263), .B1(new_n468), .B2(KEYINPUT87), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT87), .ZN(new_n470));
  AOI211_X1 g0270(.A(new_n470), .B(new_n462), .C1(new_n467), .C2(new_n465), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n453), .B(new_n455), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n206), .A2(G45), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n285), .A2(G274), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n285), .A2(G250), .A3(new_n473), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n222), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G238), .B2(G1698), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n411), .A2(new_n479), .B1(new_n283), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n373), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n355), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n472), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n462), .ZN(new_n486));
  AND4_X1   g0286(.A1(new_n207), .A2(new_n409), .A3(new_n410), .A4(new_n296), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n464), .B1(new_n487), .B2(G68), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n466), .A2(KEYINPUT86), .A3(new_n215), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n470), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n263), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n452), .A2(G87), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n482), .A2(new_n360), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G200), .B2(new_n482), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n455), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n485), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT88), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT88), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n485), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n466), .A2(new_n503), .A3(new_n217), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n207), .A2(G87), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n301), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n207), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n223), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n283), .A2(new_n480), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n207), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT24), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n463), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n506), .A4(new_n511), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n263), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT25), .ZN(new_n519));
  AOI211_X1 g0319(.A(G107), .B(new_n271), .C1(KEYINPUT92), .C2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(new_n223), .B2(new_n451), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n218), .A2(new_n302), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G257), .B2(new_n302), .ZN(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n411), .A2(new_n528), .B1(new_n283), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT5), .B(G41), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n373), .B1(new_n474), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n530), .A2(new_n373), .B1(new_n532), .B2(G264), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n531), .A2(new_n285), .A3(G274), .A4(new_n474), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(G190), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n518), .A2(new_n526), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n342), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n533), .A2(new_n355), .A3(new_n534), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n328), .B1(new_n513), .B2(new_n516), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n525), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n538), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n539), .B1(new_n538), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n480), .B1(new_n206), .B2(G33), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n273), .A2(new_n275), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n272), .A2(new_n480), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(new_n283), .B2(G97), .ZN(new_n552));
  INV_X1    g0352(.A(G283), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n283), .B2(new_n553), .ZN(new_n554));
  AOI221_X4 g0354(.A(KEYINPUT89), .B1(new_n480), .B2(G20), .C1(new_n262), .C2(new_n235), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT89), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n480), .A2(G20), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n263), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n554), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT20), .B(new_n554), .C1(new_n555), .C2(new_n558), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n551), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n224), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G257), .B2(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n463), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n301), .A2(G303), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n285), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n531), .A2(new_n474), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(G270), .A3(new_n285), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n534), .ZN(new_n572));
  OAI21_X1  g0372(.A(G169), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n547), .B1(new_n563), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n549), .A2(new_n550), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n263), .A2(new_n557), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT89), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n263), .A2(new_n556), .A3(new_n557), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT20), .B1(new_n579), .B2(new_n554), .ZN(new_n580));
  INV_X1    g0380(.A(new_n562), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n571), .A2(new_n534), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n568), .B1(new_n411), .B2(new_n565), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n373), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n342), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(KEYINPUT21), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n574), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(G179), .A3(new_n585), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT90), .B1(new_n563), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT90), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n569), .A2(new_n572), .A3(new_n355), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n582), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT91), .ZN(new_n596));
  OAI21_X1  g0396(.A(G200), .B1(new_n569), .B2(new_n572), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n563), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n563), .B2(new_n597), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n569), .A2(new_n360), .A3(new_n572), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n302), .A2(G244), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n411), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n302), .A2(KEYINPUT4), .A3(G244), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n218), .B2(new_n302), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n305), .B1(G33), .B2(G283), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n373), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n570), .A2(G257), .A3(new_n285), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n534), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT85), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n613), .A3(new_n534), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n272), .A2(new_n456), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n451), .B2(new_n456), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT6), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n456), .A2(new_n223), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n458), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n623), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n395), .A2(new_n398), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G107), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n618), .B1(new_n627), .B2(new_n263), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n285), .B1(new_n604), .B2(new_n607), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n611), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G190), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n616), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n627), .A2(new_n263), .ZN(new_n633));
  INV_X1    g0433(.A(new_n618), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n342), .B1(new_n629), .B2(new_n611), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n609), .A2(new_n612), .A3(new_n355), .A4(new_n614), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n595), .A2(new_n601), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n450), .A2(new_n502), .A3(new_n546), .A4(new_n640), .ZN(G372));
  INV_X1    g0441(.A(new_n498), .ZN(new_n642));
  INV_X1    g0442(.A(new_n638), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT26), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n638), .B1(new_n499), .B2(new_n501), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n594), .A2(new_n543), .A3(new_n574), .A4(new_n587), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT94), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n632), .A2(new_n638), .A3(new_n538), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT94), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n588), .A2(new_n650), .A3(new_n543), .A4(new_n594), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(new_n642), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n485), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n450), .B1(new_n646), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT95), .ZN(new_n655));
  INV_X1    g0455(.A(new_n357), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n326), .A2(new_n282), .B1(new_n319), .B2(new_n386), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n430), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n435), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n448), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n656), .B1(new_n661), .B2(new_n368), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(G369));
  NAND3_X1  g0463(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n542), .B2(new_n525), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n546), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT96), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n546), .A2(KEYINPUT96), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n669), .B1(new_n588), .B2(new_n594), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n543), .ZN(new_n677));
  INV_X1    g0477(.A(new_n669), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT97), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n676), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n595), .A2(new_n601), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n582), .A2(new_n669), .ZN(new_n686));
  MUX2_X1   g0486(.A(new_n595), .B(new_n685), .S(new_n686), .Z(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n673), .A2(new_n674), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n677), .A2(new_n669), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(G399));
  NAND2_X1  g0493(.A1(new_n210), .A2(new_n284), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n459), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n234), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT26), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n645), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n642), .A2(new_n649), .A3(new_n647), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT26), .B1(new_n498), .B2(new_n638), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n485), .A3(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT29), .B(new_n678), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n652), .A2(new_n485), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n485), .A2(new_n497), .A3(new_n500), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n500), .B1(new_n485), .B2(new_n497), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT26), .B(new_n643), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n700), .B1(new_n498), .B2(new_n638), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n669), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n706), .B1(new_n713), .B2(KEYINPUT29), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n592), .A2(new_n482), .A3(new_n533), .A4(new_n630), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n482), .A2(new_n533), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n589), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(new_n630), .ZN(new_n721));
  AOI211_X1 g0521(.A(G179), .B(new_n482), .C1(new_n585), .C2(new_n583), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n615), .A2(new_n536), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n717), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n724), .A2(new_n725), .A3(new_n678), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n722), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n720), .B1(new_n719), .B2(new_n630), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT98), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT98), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n733), .A3(new_n669), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n726), .B1(new_n734), .B2(new_n725), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n502), .A2(new_n640), .A3(new_n546), .A4(new_n678), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n715), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n714), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n699), .B1(new_n740), .B2(G1), .ZN(G364));
  INV_X1    g0541(.A(new_n688), .ZN(new_n742));
  INV_X1    g0542(.A(new_n694), .ZN(new_n743));
  INV_X1    g0543(.A(G13), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n206), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G330), .B2(new_n687), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n235), .B1(G20), .B2(new_n342), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n360), .A2(G179), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n207), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(new_n355), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G311), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n754), .A2(new_n529), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n755), .A2(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n360), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n759), .B1(G326), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT99), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n207), .A2(G179), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n360), .A3(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n756), .ZN(new_n766));
  INV_X1    g0566(.A(G329), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n765), .A2(new_n553), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT100), .Z(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n755), .A2(G190), .A3(new_n389), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n301), .B1(new_n770), .B2(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n760), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(KEYINPUT101), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT101), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n763), .A2(new_n769), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n761), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT32), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n766), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n783), .A2(new_n202), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G68), .B2(new_n775), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n305), .B1(new_n757), .B2(new_n221), .ZN(new_n789));
  INV_X1    g0589(.A(new_n773), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G58), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n754), .A2(new_n456), .ZN(new_n792));
  INV_X1    g0592(.A(new_n770), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(G87), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n765), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n784), .A2(new_n786), .B1(new_n795), .B2(G107), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n788), .A2(new_n791), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n752), .B1(new_n782), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n210), .A2(new_n305), .ZN(new_n799));
  INV_X1    g0599(.A(G355), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n800), .B1(G116), .B2(new_n210), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n256), .A2(G45), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n210), .A2(new_n411), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n234), .B2(new_n286), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n751), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n748), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n808), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n687), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n750), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  INV_X1    g0616(.A(new_n757), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n775), .A2(G283), .B1(new_n817), .B2(G116), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT102), .Z(new_n819));
  OAI21_X1  g0619(.A(new_n301), .B1(new_n773), .B2(new_n529), .ZN(new_n820));
  INV_X1    g0620(.A(new_n766), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(G311), .B2(new_n821), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n217), .A2(new_n765), .B1(new_n770), .B2(new_n223), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n792), .B(new_n823), .C1(G303), .C2(new_n761), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n819), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT103), .B(G143), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n790), .A2(new_n827), .B1(new_n817), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n776), .B2(new_n829), .C1(new_n830), .C2(new_n783), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n411), .B1(new_n821), .B2(G132), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n795), .A2(G68), .ZN(new_n835));
  INV_X1    g0635(.A(new_n754), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G58), .B1(new_n793), .B2(G50), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n831), .A2(new_n832), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n825), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n751), .ZN(new_n841));
  INV_X1    g0641(.A(new_n748), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n751), .A2(new_n806), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n221), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT104), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n385), .B2(new_n678), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n390), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n385), .A2(new_n845), .A3(new_n678), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n387), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n386), .A2(new_n678), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n841), .B(new_n844), .C1(new_n852), .C2(new_n807), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n713), .A2(new_n852), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT105), .B1(new_n713), .B2(new_n852), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n738), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n842), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n738), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n853), .B1(new_n861), .B2(new_n862), .ZN(G384));
  OAI211_X1 g0663(.A(G116), .B(new_n236), .C1(new_n623), .C2(KEYINPUT35), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(KEYINPUT106), .B1(KEYINPUT35), .B2(new_n623), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT106), .B2(new_n864), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n697), .A2(new_n221), .A3(new_n400), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n215), .A2(G50), .ZN(new_n869));
  OAI211_X1 g0669(.A(G1), .B(new_n744), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT107), .Z(new_n872));
  OAI21_X1  g0672(.A(new_n669), .B1(new_n724), .B2(new_n732), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n730), .A2(KEYINPUT98), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n725), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n731), .A2(new_n733), .A3(KEYINPUT31), .A4(new_n669), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n736), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n326), .A2(new_n282), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n282), .A2(new_n669), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n319), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n282), .B(new_n669), .C1(new_n320), .C2(new_n326), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n851), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n885), .A2(new_n393), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n415), .A2(new_n263), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n419), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n667), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n445), .A2(new_n447), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n660), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n442), .A2(new_n888), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n417), .A2(new_n419), .A3(new_n428), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n443), .A2(new_n889), .ZN(new_n898));
  XNOR2_X1  g0698(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n444), .A2(new_n898), .A3(new_n895), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n884), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n444), .A2(new_n898), .A3(new_n895), .ZN(new_n909));
  INV_X1    g0709(.A(new_n899), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT110), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n900), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n909), .A2(new_n912), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n898), .B1(new_n437), .B2(new_n448), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n903), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n883), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n908), .B1(new_n918), .B2(new_n907), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT112), .Z(new_n920));
  AND2_X1   g0720(.A1(new_n450), .A2(new_n877), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n715), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n921), .B2(new_n920), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n678), .B(new_n852), .C1(new_n646), .C2(new_n653), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n850), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n880), .A2(new_n881), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(new_n906), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n892), .A2(new_n667), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n878), .A2(new_n669), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n893), .B2(new_n901), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT39), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT109), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n917), .A2(new_n935), .A3(new_n905), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(KEYINPUT39), .C1(new_n931), .C2(new_n932), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n929), .B1(new_n930), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n706), .B(new_n450), .C1(new_n713), .C2(KEYINPUT29), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n662), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT111), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n941), .B(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n923), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n947), .B1(new_n206), .B2(new_n745), .C1(new_n945), .C2(new_n923), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n872), .B1(new_n948), .B2(new_n949), .ZN(G367));
  OAI211_X1 g0750(.A(new_n632), .B(new_n638), .C1(new_n628), .C2(new_n678), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n638), .B2(new_n678), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n691), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT115), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n493), .A2(new_n455), .A3(new_n494), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n669), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT114), .Z(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(new_n485), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n642), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n954), .B(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n673), .A2(new_n674), .A3(new_n675), .A4(new_n952), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n638), .B1(new_n951), .B2(new_n543), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(KEYINPUT42), .B1(new_n678), .B2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n964), .A2(new_n966), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n962), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n684), .A2(new_n952), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT45), .Z(new_n970));
  NOR2_X1   g0770(.A1(new_n684), .A2(new_n952), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n691), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n689), .A2(new_n690), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n676), .B1(new_n975), .B2(new_n675), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n688), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n739), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n970), .A2(new_n692), .A3(new_n972), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n740), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n694), .B(KEYINPUT41), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n746), .B(KEYINPUT116), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n968), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n809), .B1(new_n210), .B2(new_n454), .C1(new_n246), .C2(new_n803), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n842), .B1(new_n987), .B2(KEYINPUT117), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(KEYINPUT117), .B2(new_n987), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n790), .A2(G150), .B1(new_n821), .B2(G137), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n305), .C1(new_n202), .C2(new_n757), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n795), .A2(G77), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n253), .B2(new_n770), .C1(new_n776), .C2(new_n785), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n783), .A2(new_n826), .B1(new_n215), .B2(new_n754), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT119), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n783), .A2(new_n758), .B1(new_n223), .B2(new_n754), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n463), .B(new_n997), .C1(G97), .C2(new_n795), .ZN(new_n998));
  INV_X1    g0798(.A(G317), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n773), .A2(new_n771), .B1(new_n766), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G283), .B2(new_n817), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT118), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n770), .A2(new_n480), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n776), .A2(new_n529), .B1(KEYINPUT46), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT46), .B2(new_n1003), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n998), .B(new_n1001), .C1(new_n1002), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT118), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n996), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n989), .B1(new_n1010), .B2(new_n751), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n960), .B2(new_n813), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n986), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n977), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n985), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n689), .A2(new_n690), .A3(new_n808), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n799), .A2(new_n695), .B1(G107), .B2(new_n210), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n243), .A2(new_n286), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n695), .ZN(new_n1021));
  AOI211_X1 g0821(.A(G45), .B(new_n1021), .C1(G68), .C2(G77), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n332), .A2(G50), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n803), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1019), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n748), .B1(new_n1026), .B2(new_n810), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n770), .A2(new_n221), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n454), .A2(new_n754), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G159), .C2(new_n761), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n333), .A2(new_n775), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n773), .A2(new_n202), .B1(new_n766), .B2(new_n829), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G68), .B2(new_n817), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n411), .B1(new_n795), .B2(G97), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n463), .B1(G326), .B2(new_n821), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n754), .A2(new_n553), .B1(new_n770), .B2(new_n529), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n790), .A2(G317), .B1(new_n817), .B2(G303), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n776), .B2(new_n758), .C1(new_n772), .C2(new_n783), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1036), .B1(new_n480), .B2(new_n765), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1035), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1027), .B1(new_n1046), .B2(new_n751), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n978), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n743), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1016), .A2(new_n740), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  INV_X1    g0852(.A(new_n979), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n692), .B1(new_n970), .B2(new_n972), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n980), .A3(new_n743), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n251), .A2(new_n210), .A3(new_n411), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n809), .B1(new_n456), .B2(new_n210), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n748), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n952), .A2(new_n813), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n776), .A2(new_n771), .B1(new_n480), .B2(new_n754), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n301), .B1(new_n766), .B2(new_n772), .C1(new_n529), .C2(new_n757), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n223), .A2(new_n765), .B1(new_n770), .B2(new_n553), .ZN(new_n1063));
  OR3_X1    g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G317), .A2(new_n761), .B1(new_n790), .B2(G311), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n761), .B1(new_n790), .B2(G159), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n754), .A2(new_n221), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G50), .B2(new_n775), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n757), .A2(new_n332), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n821), .B2(new_n827), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n793), .A2(G68), .B1(new_n795), .B2(G87), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n463), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1064), .A2(new_n1066), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1059), .B(new_n1060), .C1(new_n751), .C2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n1017), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1056), .A2(new_n1078), .ZN(G390));
  AND3_X1   g0879(.A1(new_n737), .A2(KEYINPUT121), .A3(new_n882), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT121), .B1(new_n737), .B2(new_n882), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n917), .A2(new_n905), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n930), .B(KEYINPUT120), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n850), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n705), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n669), .B1(new_n1086), .B2(new_n701), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1087), .B2(new_n849), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n926), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1083), .B(new_n1084), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n930), .B1(new_n925), .B2(new_n926), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1082), .B(new_n1090), .C1(new_n939), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n877), .A2(new_n882), .A3(G330), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n938), .A2(new_n936), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n930), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1085), .B1(new_n713), .B2(new_n852), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n1089), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1099), .A3(new_n934), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1095), .B1(new_n1100), .B2(new_n1090), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n450), .A2(G330), .A3(new_n877), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n942), .A2(new_n1102), .A3(new_n662), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT122), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n942), .A2(new_n1102), .A3(new_n662), .A4(KEYINPUT122), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n926), .B1(new_n737), .B2(new_n852), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n925), .B1(new_n1108), .B2(new_n1094), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n877), .A2(G330), .A3(new_n852), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1089), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1088), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1093), .A2(new_n1101), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1114), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1090), .B1(new_n939), .B2(new_n1091), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1094), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1092), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1120), .A3(new_n743), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1096), .A2(new_n806), .A3(new_n934), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n843), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n748), .B1(new_n333), .B2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n836), .A2(G159), .B1(new_n817), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n830), .B2(new_n776), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT123), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n793), .A2(G150), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  INV_X1    g0933(.A(G132), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n305), .B1(new_n766), .B2(new_n1133), .C1(new_n773), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(G128), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n783), .A2(new_n1136), .B1(new_n765), .B2(new_n202), .ZN(new_n1137));
  OR3_X1    g0937(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1069), .B1(G283), .B2(new_n761), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n223), .B2(new_n776), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n773), .A2(new_n480), .B1(new_n766), .B2(new_n529), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n305), .B(new_n1141), .C1(G97), .C2(new_n817), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n793), .A2(G87), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n835), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1130), .A2(new_n1138), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1125), .B1(new_n1145), .B2(new_n751), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1122), .A2(new_n1017), .B1(new_n1123), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1121), .A2(new_n1147), .ZN(G378));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n907), .B1(new_n1083), .B2(new_n884), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n877), .A2(new_n882), .A3(new_n907), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n905), .B2(new_n904), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n368), .A2(new_n357), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n341), .A2(new_n667), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1156), .B(new_n1157), .Z(new_n1160));
  NAND3_X1  g0960(.A1(new_n919), .A2(new_n1160), .A3(G330), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n941), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n940), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1149), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1120), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1120), .A2(new_n1166), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n743), .C1(KEYINPUT57), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n842), .B1(new_n202), .B2(new_n843), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1133), .A2(new_n783), .B1(new_n776), .B2(new_n1134), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n790), .A2(G128), .B1(new_n817), .B2(G137), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n770), .B2(new_n1126), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G150), .C2(new_n836), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n795), .A2(G159), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n821), .C2(G124), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n790), .A2(G107), .B1(new_n821), .B2(G283), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n454), .B2(new_n757), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1028), .B(new_n1183), .C1(G68), .C2(new_n836), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n783), .A2(new_n480), .B1(new_n765), .B2(new_n253), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G97), .B2(new_n775), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1184), .A2(new_n284), .A3(new_n411), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT58), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G50), .B1(new_n283), .B2(new_n284), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n463), .B2(G41), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n1181), .A2(new_n1189), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1171), .B1(new_n752), .B2(new_n1193), .C1(new_n1160), .C2(new_n807), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n1017), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1170), .A2(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1089), .A2(new_n806), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n480), .A2(new_n776), .B1(new_n783), .B2(new_n529), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G97), .B2(new_n793), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1029), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n773), .A2(new_n553), .B1(new_n757), .B2(new_n223), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n305), .B(new_n1203), .C1(G303), .C2(new_n821), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n992), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n757), .A2(new_n829), .B1(new_n766), .B2(new_n1136), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G137), .B2(new_n790), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G50), .A2(new_n836), .B1(new_n775), .B2(new_n1127), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n761), .A2(G132), .B1(new_n793), .B2(G159), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n411), .B1(new_n795), .B2(G58), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n752), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n842), .B(new_n1212), .C1(new_n215), .C2(new_n843), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1114), .A2(new_n1017), .B1(new_n1199), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1166), .A2(new_n1114), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n983), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1166), .A2(new_n1114), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(G381));
  OR4_X1    g1018(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(G387), .A3(G381), .ZN(new_n1220));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1220), .A2(new_n1221), .A3(new_n1170), .A4(new_n1197), .ZN(G407));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n668), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  XNOR2_X1  g1024(.A(G393), .B(new_n815), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G390), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1225), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1056), .A3(new_n1078), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1014), .A2(new_n1226), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1228), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1227), .B1(new_n1056), .B2(new_n1078), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1230), .A2(new_n1231), .B1(new_n986), .B2(new_n1013), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n668), .A2(G213), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1107), .B1(new_n1122), .B2(new_n1117), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n940), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n939), .A2(new_n930), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n929), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1159), .A2(new_n1161), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n743), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1196), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G378), .B(new_n1197), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1170), .A2(KEYINPUT124), .A3(G378), .A4(new_n1197), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1169), .A2(new_n983), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1197), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1221), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1235), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1235), .A2(G2897), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1217), .B1(KEYINPUT60), .B2(new_n1215), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1107), .A2(new_n1115), .A3(KEYINPUT60), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n743), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1214), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G384), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1253), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1253), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1234), .B1(new_n1252), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1252), .B2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1246), .A2(new_n1247), .B1(new_n1221), .B2(new_n1250), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(new_n1267), .A3(new_n1235), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1266), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1233), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1233), .B1(KEYINPUT63), .B2(new_n1272), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1263), .B(new_n1262), .C1(new_n1271), .C2(new_n1235), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1234), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT125), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1233), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1273), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1277), .B(new_n1234), .C1(new_n1272), .C2(new_n1266), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1272), .A2(KEYINPUT63), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1265), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1233), .A4(new_n1276), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1280), .A2(new_n1289), .ZN(G405));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G375), .A2(new_n1221), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(KEYINPUT126), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1293), .B2(new_n1248), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1291), .A3(new_n1248), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1267), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1296), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1298), .A2(new_n1268), .A3(new_n1294), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1281), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1268), .B1(new_n1298), .B2(new_n1294), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1295), .A2(new_n1267), .A3(new_n1296), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1233), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(G402));
endmodule


