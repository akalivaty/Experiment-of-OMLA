//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT69), .ZN(new_n458));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(G567), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(KEYINPUT69), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n464), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT70), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT72), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n465), .A2(new_n466), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(G136), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n481), .B2(new_n464), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n465), .B2(new_n466), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n499), .B(new_n502), .C1(new_n466), .C2(new_n465), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(G166));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n516));
  AND3_X1   g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n505), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n521), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n534), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AND2_X1   g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n522), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT75), .B(G90), .Z(new_n546));
  AOI22_X1  g121(.A1(G651), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n538), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n534), .A2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n542), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT76), .B(G81), .Z(new_n554));
  AOI22_X1  g129(.A1(G651), .A2(new_n553), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT77), .B1(new_n509), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n531), .A2(new_n565), .A3(G53), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n564), .A2(KEYINPUT9), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g143(.A(KEYINPUT77), .B(new_n568), .C1(new_n509), .C2(new_n563), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n542), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n545), .A2(G91), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(G166), .A2(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(new_n511), .B2(new_n514), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G303));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n513), .B1(new_n542), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(G87), .B2(new_n545), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n531), .A2(KEYINPUT79), .A3(G49), .ZN(new_n585));
  OAI211_X1 g160(.A(G49), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n584), .A2(new_n589), .ZN(G288));
  OAI21_X1  g165(.A(G61), .B1(new_n540), .B2(new_n541), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI211_X1 g167(.A(KEYINPUT80), .B(new_n513), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n507), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT80), .B1(new_n598), .B2(new_n513), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n542), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G85), .B2(new_n545), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n534), .A2(G47), .B1(new_n604), .B2(KEYINPUT81), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n534), .A2(G54), .ZN(new_n610));
  INV_X1    g185(.A(G79), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n611), .A2(new_n528), .A3(KEYINPUT82), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT82), .B1(new_n611), .B2(new_n528), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n542), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G651), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n545), .A2(KEYINPUT10), .A3(G92), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n507), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n610), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n576), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(G868), .B2(new_n576), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(G148));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n556), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n622), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n488), .A2(G123), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(G111), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G2105), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n482), .B2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n486), .A2(new_n468), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT13), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(G2100), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n648), .B2(new_n647), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n644), .A2(new_n645), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT85), .B(G2438), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n661), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT87), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n685), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n685), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT89), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n717), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n709), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n709), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G1971), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  INV_X1    g300(.A(G305), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G16), .ZN(new_n727));
  OR2_X1    g302(.A1(G6), .A2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT32), .B(G1981), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT88), .ZN(new_n732));
  OAI21_X1  g307(.A(KEYINPUT88), .B1(new_n730), .B2(new_n731), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n724), .A2(new_n725), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT34), .B1(new_n735), .B2(new_n723), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G24), .ZN(new_n737));
  INV_X1    g312(.A(G290), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n709), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1986), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n488), .A2(G119), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n482), .A2(G131), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n464), .A2(G107), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  MUX2_X1   g320(.A(G25), .B(new_n745), .S(G29), .Z(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n746), .B(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n740), .A2(KEYINPUT90), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n734), .A2(new_n736), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n488), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n468), .A2(G105), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT97), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n482), .A2(G141), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n755), .A2(new_n757), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n754), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n754), .A2(G32), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT27), .B(G1996), .Z(new_n769));
  OAI21_X1  g344(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n754), .A2(G33), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n486), .A2(G127), .ZN(new_n775));
  AND2_X1   g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  OAI21_X1  g351(.A(G2105), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT93), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(KEYINPUT93), .B(G2105), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  NAND2_X1  g356(.A1(G103), .A2(G2104), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n482), .A2(G139), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n779), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT94), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT95), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n774), .B1(new_n788), .B2(G29), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n773), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n557), .A2(new_n709), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n709), .B2(G19), .ZN(new_n793));
  INV_X1    g368(.A(G1341), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n754), .A2(G27), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT104), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n501), .A2(new_n503), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n492), .A2(new_n496), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n754), .B1(new_n483), .B2(new_n489), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n754), .A2(G35), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n804), .A2(KEYINPUT29), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G2090), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT29), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n709), .A2(G5), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G171), .B2(new_n709), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n793), .A2(new_n794), .B1(new_n811), .B2(G1961), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n803), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(G160), .A2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT24), .B(G34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n754), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT96), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2084), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n754), .A2(G26), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n488), .A2(G128), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n825));
  INV_X1    g400(.A(G116), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G2105), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n482), .B2(G140), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n823), .B1(new_n829), .B2(G29), .ZN(new_n830));
  INV_X1    g405(.A(G2067), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G4), .A2(G16), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT91), .Z(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n622), .B2(new_n709), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1348), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n791), .A2(new_n813), .A3(new_n833), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n790), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n643), .A2(new_n754), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT101), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n709), .A2(G21), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G286), .B2(G16), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT100), .B(G1966), .Z(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G1961), .B2(new_n811), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT31), .B(G11), .ZN(new_n847));
  INV_X1    g422(.A(G28), .ZN(new_n848));
  AOI21_X1  g423(.A(G29), .B1(new_n848), .B2(KEYINPUT30), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT102), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(KEYINPUT30), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n849), .A2(KEYINPUT102), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n843), .B2(new_n844), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT103), .B1(new_n841), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n840), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(new_n859), .A3(new_n854), .A4(new_n846), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n709), .A2(G20), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT23), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n576), .B2(new_n709), .ZN(new_n864));
  INV_X1    g439(.A(G1956), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n806), .A2(new_n808), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n807), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n861), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n734), .A2(KEYINPUT36), .A3(new_n736), .A4(new_n750), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n753), .A2(new_n839), .A3(new_n871), .A4(new_n872), .ZN(G150));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n874));
  XNOR2_X1  g449(.A(G150), .B(new_n874), .ZN(G311));
  NAND2_X1  g450(.A1(new_n534), .A2(G55), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n877));
  NAND2_X1  g452(.A1(G80), .A2(G543), .ZN(new_n878));
  INV_X1    g453(.A(G67), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n542), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(G651), .A2(new_n880), .B1(new_n545), .B2(G93), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n877), .B1(new_n876), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n556), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(new_n881), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n556), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n623), .A2(G559), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n893));
  AOI21_X1  g468(.A(G860), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n886), .A2(KEYINPUT107), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n882), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G860), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT37), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(G145));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n901));
  INV_X1    g476(.A(new_n503), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n502), .B1(new_n486), .B2(new_n499), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n904), .B2(new_n497), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT109), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n764), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n761), .A2(new_n762), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n763), .A2(new_n764), .A3(new_n907), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n829), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n829), .B1(new_n911), .B2(new_n912), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n788), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n787), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n482), .A2(G142), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n464), .A2(G118), .ZN(new_n920));
  OAI21_X1  g495(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(G130), .B2(new_n488), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(new_n647), .Z(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(new_n745), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n918), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n916), .A2(new_n918), .A3(new_n928), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n916), .A2(new_n918), .ZN(new_n930));
  INV_X1    g505(.A(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(G160), .B(KEYINPUT108), .Z(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(G162), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(G162), .ZN(new_n936));
  INV_X1    g511(.A(new_n643), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n925), .B1(new_n916), .B2(new_n918), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n940), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n943), .B2(new_n926), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT40), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT40), .B1(new_n941), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(G395));
  NAND2_X1  g522(.A1(new_n897), .A2(new_n631), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n889), .B(new_n633), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n576), .A2(new_n622), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT111), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n576), .A2(new_n622), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n576), .A2(new_n954), .A3(new_n622), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n953), .A3(new_n958), .A4(new_n955), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n949), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n961));
  INV_X1    g536(.A(new_n955), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n954), .B1(new_n576), .B2(new_n622), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n951), .A2(KEYINPUT113), .A3(new_n955), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n952), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n951), .A2(new_n955), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n953), .A2(KEYINPUT41), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n966), .A2(KEYINPUT41), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n960), .B1(new_n949), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(G166), .B(KEYINPUT114), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n971), .A2(new_n726), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n726), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(G290), .B(G288), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n738), .A2(G288), .ZN(new_n977));
  NOR2_X1   g552(.A1(G290), .A2(new_n711), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n977), .A2(new_n978), .B1(new_n972), .B2(new_n973), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n970), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n948), .B1(new_n982), .B2(new_n631), .ZN(G295));
  OAI21_X1  g558(.A(new_n948), .B1(new_n982), .B2(new_n631), .ZN(G331));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n985));
  INV_X1    g560(.A(new_n956), .ZN(new_n986));
  NAND3_X1  g561(.A1(G286), .A2(new_n538), .A3(new_n547), .ZN(new_n987));
  NAND3_X1  g562(.A1(G301), .A2(new_n535), .A3(new_n526), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n885), .A2(new_n888), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n557), .B1(new_n896), .B2(new_n882), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n887), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n986), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n989), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n969), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n980), .ZN(new_n997));
  AOI21_X1  g572(.A(G37), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n993), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n967), .A2(new_n968), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n962), .A2(new_n961), .A3(new_n963), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT113), .B1(new_n951), .B2(new_n955), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n953), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT41), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n999), .B1(new_n1005), .B2(new_n994), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n980), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n985), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n993), .B(new_n980), .C1(new_n969), .C2(new_n995), .ZN(new_n1009));
  INV_X1    g584(.A(G37), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n994), .A2(new_n957), .A3(new_n959), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n980), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n986), .A2(KEYINPUT41), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n968), .B1(new_n964), .B2(new_n965), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n994), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1010), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1009), .A2(new_n1016), .A3(KEYINPUT43), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1008), .A2(new_n1017), .A3(KEYINPUT44), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n998), .A2(new_n985), .A3(new_n1007), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n998), .A2(KEYINPUT115), .A3(new_n1007), .A4(new_n985), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT43), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1024), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n907), .B2(G1384), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n471), .A2(new_n475), .A3(G40), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n829), .B(new_n831), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n745), .A2(new_n748), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n763), .A2(new_n764), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G1996), .ZN(new_n1035));
  INV_X1    g610(.A(G1996), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1031), .B(new_n1032), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n824), .A2(new_n831), .A3(new_n828), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1030), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1030), .A2(G1986), .A3(G290), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1041), .B(KEYINPUT48), .Z(new_n1042));
  XNOR2_X1  g617(.A(new_n745), .B(new_n747), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1031), .B(new_n1043), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n1029), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1040), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT126), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1030), .B1(new_n1034), .B2(new_n1031), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1046), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT127), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1046), .B(KEYINPUT127), .C1(new_n1055), .C2(new_n1054), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n798), .B2(new_n799), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n1064));
  INV_X1    g639(.A(G40), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(new_n470), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1062), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n597), .B2(new_n599), .ZN(new_n1069));
  INV_X1    g644(.A(new_n596), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n591), .A2(new_n592), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT80), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(G651), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT118), .B(G1981), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1070), .A2(new_n599), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT119), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n597), .A2(new_n1077), .A3(new_n599), .A4(new_n1074), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1069), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1067), .B1(new_n1079), .B2(KEYINPUT49), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1081), .B(new_n1069), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G288), .A2(G1976), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1083), .A2(new_n1084), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1067), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n578), .A2(G8), .A3(new_n580), .ZN(new_n1087));
  XOR2_X1   g662(.A(new_n1087), .B(KEYINPUT55), .Z(new_n1088));
  INV_X1    g663(.A(G1384), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n800), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1028), .B1(new_n1090), .B2(new_n1026), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n905), .A2(KEYINPUT45), .A3(new_n1089), .A4(new_n906), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1971), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(KEYINPUT116), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(new_n1089), .C1(new_n904), .C2(new_n497), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1066), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1093), .A2(KEYINPUT116), .B1(G2090), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1088), .B(G8), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1976), .B1(new_n584), .B2(new_n589), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT52), .B1(new_n1067), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n584), .A2(new_n589), .A3(G1976), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(G8), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1105), .A2(new_n1104), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(new_n1067), .C1(KEYINPUT52), .C2(new_n1101), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1085), .A2(new_n1086), .B1(new_n1100), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1087), .B(KEYINPUT55), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1098), .A2(G2090), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n1093), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G8), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1093), .A2(new_n1115), .A3(KEYINPUT120), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1111), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1110), .B(KEYINPUT121), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1119), .A2(new_n1100), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1066), .B1(new_n1063), .B2(KEYINPUT45), .ZN(new_n1124));
  NOR3_X1   g699(.A1(G164), .A2(new_n1026), .A3(G1384), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n844), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1095), .A2(new_n1097), .A3(new_n819), .A4(new_n1066), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G8), .A3(G168), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1113), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(G8), .B1(new_n1099), .B2(new_n1094), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1114), .A2(KEYINPUT122), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1111), .A2(new_n1113), .A3(new_n1129), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1112), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1123), .ZN(new_n1138));
  INV_X1    g713(.A(G2078), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1091), .A2(new_n1092), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT53), .ZN(new_n1141));
  INV_X1    g716(.A(G1961), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1140), .A2(new_n1141), .B1(new_n1142), .B2(new_n1098), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n800), .A2(KEYINPUT45), .A3(new_n1089), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1141), .A2(G2078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1091), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G301), .B(KEYINPUT54), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1092), .A2(new_n1066), .A3(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1027), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1147), .A2(new_n1148), .B1(new_n1150), .B2(new_n1143), .ZN(new_n1151));
  NAND2_X1  g726(.A1(G286), .A2(G8), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1095), .A2(new_n1066), .A3(new_n1097), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1026), .B1(G164), .B2(G1384), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(new_n1144), .A3(new_n1066), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1157), .A2(new_n819), .B1(new_n1159), .B2(new_n844), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1152), .B(new_n1156), .C1(new_n1160), .C2(new_n1062), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT51), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1162));
  OAI211_X1 g737(.A(G8), .B(new_n1162), .C1(new_n1128), .C2(G286), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1128), .A2(G8), .A3(G286), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1151), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1091), .A2(new_n1092), .A3(new_n1036), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1103), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n556), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1063), .A2(new_n831), .A3(new_n1066), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1063), .A2(KEYINPUT123), .A3(new_n1066), .A4(new_n831), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G1348), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1098), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1175), .A2(new_n1176), .B1(new_n1098), .B2(new_n1178), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n622), .B1(new_n1183), .B2(KEYINPUT60), .ZN(new_n1184));
  AND4_X1   g759(.A1(KEYINPUT60), .A2(new_n1177), .A3(new_n1179), .A4(new_n622), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1182), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT57), .B1(new_n567), .B2(new_n575), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n573), .A2(new_n574), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT57), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n564), .A2(KEYINPUT9), .A3(new_n566), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n569), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(KEYINPUT56), .B(G2072), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1091), .A2(new_n1092), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1098), .A2(new_n865), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1194), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1187), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n1193), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1203), .A2(KEYINPUT61), .A3(new_n1198), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1172), .A2(new_n1186), .A3(new_n1201), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1183), .A2(new_n622), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1200), .B1(new_n1206), .B2(new_n1198), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1166), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1165), .A2(KEYINPUT62), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1161), .A2(new_n1163), .A3(new_n1210), .A4(new_n1164), .ZN(new_n1211));
  AOI21_X1  g786(.A(G301), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1138), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1137), .A2(new_n1214), .ZN(new_n1215));
  XOR2_X1   g790(.A(G290), .B(G1986), .Z(new_n1216));
  INV_X1    g791(.A(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1029), .B1(new_n1044), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1061), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1218), .ZN(new_n1220));
  AOI211_X1 g795(.A(KEYINPUT125), .B(new_n1220), .C1(new_n1137), .C2(new_n1214), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1060), .B1(new_n1219), .B2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g797(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n706), .B2(new_n707), .ZN(new_n1225));
  INV_X1    g799(.A(new_n940), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n942), .B1(KEYINPUT110), .B2(new_n926), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1226), .B1(new_n1227), .B2(new_n929), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n1226), .A2(new_n926), .A3(new_n932), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1229), .A2(new_n1010), .ZN(new_n1230));
  OAI21_X1  g804(.A(new_n1225), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g805(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1232));
  NOR2_X1   g806(.A1(new_n1231), .A2(new_n1232), .ZN(G308));
  OAI221_X1 g807(.A(new_n1225), .B1(new_n1008), .B2(new_n1017), .C1(new_n1228), .C2(new_n1230), .ZN(G225));
endmodule


