//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(G237), .A2(G953), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(G214), .C1(KEYINPUT83), .C2(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n187), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT18), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT84), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n199), .B(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(new_n195), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(KEYINPUT18), .B2(G131), .ZN(new_n202));
  OR3_X1    g016(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(KEYINPUT17), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT86), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(G146), .A3(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n201), .A2(G131), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n214), .A2(KEYINPUT17), .A3(new_n196), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n205), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G113), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n203), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n203), .A2(new_n216), .ZN(new_n222));
  INV_X1    g036(.A(new_n219), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI211_X1 g038(.A(KEYINPUT87), .B(new_n219), .C1(new_n203), .C2(new_n216), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G475), .ZN(new_n229));
  INV_X1    g043(.A(G475), .ZN(new_n230));
  INV_X1    g044(.A(new_n220), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT19), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n199), .B1(KEYINPUT85), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(KEYINPUT85), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  OAI221_X1 g049(.A(new_n212), .B1(new_n196), .B2(new_n214), .C1(new_n235), .C2(G146), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n219), .B1(new_n203), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n230), .B(new_n227), .C1(new_n231), .C2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n203), .A2(new_n236), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n220), .B1(new_n241), .B2(new_n219), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT20), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n230), .A4(new_n227), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n229), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n189), .A2(G952), .ZN(new_n247));
  NAND2_X1  g061(.A1(G234), .A2(G237), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n249), .B(KEYINPUT91), .Z(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT21), .B(G898), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT92), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n254), .A2(G902), .A3(new_n248), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n255), .B2(G953), .ZN(new_n256));
  INV_X1    g070(.A(G478), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT15), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(G128), .A3(new_n192), .ZN(new_n261));
  XNOR2_X1  g075(.A(G128), .B(G143), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n261), .B(G134), .C1(new_n263), .C2(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G122), .ZN(new_n268));
  INV_X1    g082(.A(G122), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT88), .B1(new_n269), .B2(G116), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT88), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n267), .A3(G122), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n264), .B(new_n266), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT14), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n275), .B1(new_n278), .B2(new_n268), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n262), .B(new_n265), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n273), .B1(KEYINPUT14), .B2(new_n274), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT9), .B(G234), .Z(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(G217), .A3(new_n189), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n283), .A2(new_n285), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G902), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n259), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n289), .B(KEYINPUT90), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n258), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n246), .A2(new_n256), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G221), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n284), .B2(new_n227), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n210), .A2(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n192), .A2(G146), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(G128), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G143), .B(G146), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n304), .A2(KEYINPUT65), .A3(new_n300), .A4(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n307), .A2(G128), .B1(new_n298), .B2(new_n299), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n218), .A2(G107), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n218), .A2(G107), .ZN(new_n314));
  OAI21_X1  g128(.A(G101), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(new_n218), .B2(G107), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n274), .A3(G104), .ZN(new_n318));
  INV_X1    g132(.A(G101), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .A4(new_n312), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n310), .A2(new_n311), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n308), .B1(new_n303), .B2(new_n305), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT76), .B1(new_n324), .B2(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n304), .ZN(new_n327));
  OAI21_X1  g141(.A(G128), .B1(new_n307), .B2(KEYINPUT66), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n298), .B2(KEYINPUT1), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n306), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n321), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT64), .B1(new_n265), .B2(G137), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n265), .A2(G137), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT64), .B(new_n339), .C1(new_n265), .C2(G137), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G131), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n337), .A2(new_n187), .A3(new_n338), .A4(new_n340), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(KEYINPUT12), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT12), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n323), .A2(new_n325), .B1(new_n333), .B2(new_n321), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n304), .A2(KEYINPUT0), .A3(G128), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G128), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n304), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n316), .A2(new_n318), .A3(new_n312), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G101), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(G101), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT4), .A3(new_n320), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n332), .A2(KEYINPUT10), .A3(new_n322), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT77), .B1(new_n326), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n364), .B(KEYINPUT10), .C1(new_n323), .C2(new_n325), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n360), .B(new_n361), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n350), .B1(new_n366), .B2(new_n344), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n189), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT10), .B1(new_n323), .B2(new_n325), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT77), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(new_n348), .A3(new_n360), .A4(new_n361), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n344), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n370), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n377), .A3(G469), .ZN(new_n378));
  NAND2_X1  g192(.A1(G469), .A2(G902), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G469), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n370), .B(new_n350), .C1(new_n366), .C2(new_n344), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n381), .B(new_n227), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n297), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n333), .A2(new_n207), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n353), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n189), .A2(G224), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n387), .A2(new_n388), .B1(KEYINPUT7), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n391));
  INV_X1    g205(.A(G119), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G116), .ZN(new_n393));
  XOR2_X1   g207(.A(G116), .B(G119), .Z(new_n394));
  OAI211_X1 g208(.A(G113), .B(new_n393), .C1(new_n394), .C2(new_n391), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT2), .B(G113), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(new_n321), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G122), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n401), .B(KEYINPUT8), .Z(new_n402));
  AOI21_X1  g216(.A(KEYINPUT81), .B1(new_n397), .B2(new_n321), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n390), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n394), .B(new_n396), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n359), .A3(new_n357), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n359), .A3(KEYINPUT79), .A4(new_n357), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n398), .A3(new_n401), .A4(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT7), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n388), .A2(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n388), .A2(KEYINPUT80), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n387), .A2(new_n413), .A3(new_n389), .A4(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n405), .B(new_n411), .C1(new_n412), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n409), .A2(new_n398), .A3(new_n410), .ZN(new_n417));
  INV_X1    g231(.A(new_n401), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT6), .A3(new_n411), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n387), .A2(new_n413), .A3(new_n414), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(G224), .A3(new_n189), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n415), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(new_n424), .A3(new_n418), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n416), .A2(new_n426), .A3(new_n227), .ZN(new_n427));
  OAI21_X1  g241(.A(G210), .B1(G237), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n416), .A2(new_n426), .A3(new_n227), .A4(new_n428), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT78), .Z(new_n434));
  AND2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n295), .A2(new_n386), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n338), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n265), .A2(G137), .ZN(new_n438));
  OAI21_X1  g252(.A(G131), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n343), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n306), .B2(new_n331), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n353), .B1(new_n342), .B2(new_n343), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n441), .A2(new_n442), .A3(new_n406), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT28), .ZN(new_n444));
  INV_X1    g258(.A(new_n406), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n344), .A2(new_n354), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n343), .A2(new_n439), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n332), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT28), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n194), .A2(G210), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n319), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n444), .A2(new_n450), .A3(KEYINPUT29), .A4(new_n455), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n456), .A2(KEYINPUT69), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n456), .B2(KEYINPUT69), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n441), .C2(new_n442), .ZN(new_n459));
  OR2_X1    g273(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n446), .A2(new_n448), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n406), .ZN(new_n464));
  INV_X1    g278(.A(new_n443), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(new_n455), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n444), .A2(new_n450), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n454), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n457), .B(new_n458), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n445), .B1(new_n459), .B2(new_n462), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n474), .A2(new_n443), .A3(new_n454), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n475), .A2(new_n476), .B1(new_n470), .B2(new_n454), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT68), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n464), .A2(new_n465), .A3(new_n455), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT31), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT32), .ZN(new_n483));
  NOR2_X1   g297(.A1(G472), .A2(G902), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n199), .A2(new_n210), .ZN(new_n489));
  XOR2_X1   g303(.A(G119), .B(G128), .Z(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT71), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT24), .B(G110), .Z(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n392), .A2(G128), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n496));
  INV_X1    g310(.A(G128), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n495), .B(new_n496), .C1(G119), .C2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n212), .B(new_n489), .C1(new_n493), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n491), .A2(new_n492), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(G110), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n213), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT22), .B(G137), .ZN(new_n505));
  INV_X1    g319(.A(G234), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n296), .A2(new_n506), .A3(G953), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n505), .B(new_n507), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(new_n503), .A3(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n227), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT72), .B1(new_n514), .B2(KEYINPUT73), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(KEYINPUT73), .B2(KEYINPUT25), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT25), .B1(KEYINPUT72), .B2(KEYINPUT73), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G217), .B1(new_n506), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(G902), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n523), .B(KEYINPUT74), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n510), .A2(new_n511), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n473), .C1(new_n485), .C2(new_n486), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n488), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n488), .A2(new_n526), .A3(new_n531), .A4(new_n528), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n436), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n319), .ZN(G3));
  INV_X1    g348(.A(new_n433), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n430), .B2(new_n431), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n256), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n289), .A2(new_n257), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n286), .B2(new_n287), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n542), .A2(KEYINPUT94), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n288), .A2(KEYINPUT33), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(KEYINPUT94), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n540), .B1(new_n546), .B2(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n257), .A2(new_n227), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n538), .A2(new_n246), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n522), .A2(new_n525), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n482), .A2(new_n484), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n482), .B2(new_n227), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n553), .A2(new_n560), .A3(new_n386), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT34), .B(G104), .Z(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(G6));
  XNOR2_X1  g377(.A(new_n238), .B(new_n239), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n564), .A2(new_n229), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n538), .A2(new_n565), .A3(new_n294), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n386), .A3(new_n560), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G107), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT95), .B(KEYINPUT35), .Z(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G9));
  XNOR2_X1  g384(.A(new_n504), .B(KEYINPUT96), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n509), .A2(KEYINPUT36), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n524), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n519), .B2(new_n521), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n436), .A2(new_n559), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT37), .B(G110), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G12));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n580));
  INV_X1    g394(.A(new_n576), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n488), .A2(new_n528), .A3(new_n386), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(new_n537), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n189), .A2(G900), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G902), .A3(new_n248), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT97), .Z(new_n586));
  NAND2_X1  g400(.A1(new_n250), .A2(new_n586), .ZN(new_n587));
  AND4_X1   g401(.A1(new_n229), .A2(new_n564), .A3(new_n294), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n580), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n582), .A2(KEYINPUT98), .A3(new_n590), .A4(new_n537), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n497), .ZN(G30));
  XNOR2_X1  g407(.A(new_n432), .B(KEYINPUT38), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n246), .A2(new_n294), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n433), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n485), .A2(new_n486), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n467), .A2(new_n454), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n443), .A2(new_n449), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n227), .B1(new_n600), .B2(new_n455), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT99), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n587), .B(KEYINPUT39), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n386), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT40), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(KEYINPUT40), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n576), .ZN(new_n609));
  OR4_X1    g423(.A1(new_n596), .A2(new_n604), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G143), .ZN(G45));
  AOI22_X1  g425(.A1(new_n228), .A2(G475), .B1(new_n240), .B2(new_n244), .ZN(new_n612));
  INV_X1    g426(.A(new_n587), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n612), .A2(new_n550), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n583), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G146), .ZN(G48));
  AND3_X1   g430(.A1(new_n488), .A2(new_n526), .A3(new_n528), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n227), .B1(new_n382), .B2(new_n384), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G469), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n385), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n297), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n617), .A2(KEYINPUT100), .A3(new_n553), .A4(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n488), .A2(new_n526), .A3(new_n621), .A4(new_n528), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(new_n552), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT41), .B(G113), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G15));
  INV_X1    g442(.A(new_n624), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n566), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G116), .ZN(G18));
  INV_X1    g445(.A(new_n297), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n632), .A2(new_n619), .A3(new_n385), .A4(new_n536), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n488), .A2(new_n633), .A3(new_n528), .A4(new_n581), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n295), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G119), .ZN(G21));
  XNOR2_X1  g450(.A(new_n484), .B(KEYINPUT101), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n479), .A2(KEYINPUT31), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n477), .B2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n554), .A2(new_n558), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n538), .A3(new_n595), .A4(new_n621), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G122), .ZN(G24));
  NOR3_X1   g456(.A1(new_n576), .A2(new_n558), .A3(new_n639), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n614), .A3(new_n633), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G125), .ZN(G27));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n646));
  INV_X1    g460(.A(new_n385), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n378), .A2(new_n379), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT102), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n385), .A2(new_n650), .A3(new_n379), .A4(new_n378), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n632), .A3(new_n614), .A4(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n646), .B1(new_n655), .B2(new_n529), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n297), .B(new_n653), .C1(new_n649), .C2(new_n651), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n554), .B1(new_n597), .B2(new_n473), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(KEYINPUT42), .A3(new_n614), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n656), .B2(new_n659), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n187), .ZN(G33));
  NAND4_X1  g478(.A1(new_n488), .A2(new_n526), .A3(new_n588), .A4(new_n528), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n657), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n652), .A2(new_n632), .A3(new_n654), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT104), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G134), .ZN(G36));
  NAND2_X1  g486(.A1(new_n551), .A2(new_n612), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT43), .Z(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n559), .A3(new_n581), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n653), .B1(new_n675), .B2(KEYINPUT44), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n372), .A2(new_n377), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G469), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT46), .B1(new_n679), .B2(new_n379), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n647), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n679), .A2(KEYINPUT46), .A3(new_n379), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n297), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(new_n605), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n676), .B(new_n684), .C1(KEYINPUT44), .C2(new_n675), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G137), .ZN(G39));
  XNOR2_X1  g500(.A(new_n683), .B(KEYINPUT47), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n488), .A2(new_n528), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n554), .A3(new_n614), .A4(new_n654), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT105), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT106), .B(G140), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G42));
  NOR4_X1   g507(.A1(new_n620), .A2(new_n250), .A3(new_n297), .A4(new_n653), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n674), .A2(new_n658), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT48), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n551), .A2(new_n246), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n604), .A2(new_n526), .A3(new_n694), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n696), .B(new_n247), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n674), .A2(new_n251), .A3(new_n640), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n700), .A2(new_n621), .ZN(new_n701));
  INV_X1    g515(.A(new_n594), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n535), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT50), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n698), .A2(new_n246), .A3(new_n551), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(KEYINPUT51), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n674), .A2(new_n643), .A3(new_n694), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n620), .A2(new_n632), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n654), .B(new_n700), .C1(new_n687), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n706), .A3(KEYINPUT51), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n706), .A2(KEYINPUT51), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n714), .A3(new_n709), .A4(new_n711), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n699), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n650), .B1(new_n380), .B2(new_n385), .ZN(new_n717));
  INV_X1    g531(.A(new_n651), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n632), .B(new_n576), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT110), .B1(new_n719), .B2(new_n613), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n595), .A2(new_n432), .A3(new_n433), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n297), .B1(new_n649), .B2(new_n651), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n576), .A4(new_n587), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n603), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n723), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n726), .A2(new_n603), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n724), .A2(new_n576), .A3(new_n587), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n721), .B1(new_n731), .B2(KEYINPUT110), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT111), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n615), .B(new_n644), .C1(new_n589), .C2(new_n591), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n615), .A2(new_n644), .ZN(new_n738));
  INV_X1    g552(.A(new_n589), .ZN(new_n739));
  INV_X1    g553(.A(new_n591), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n728), .B1(new_n723), .B2(new_n727), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n730), .A2(KEYINPUT111), .A3(new_n732), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n737), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n657), .A2(new_n614), .A3(new_n643), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n565), .A2(new_n587), .A3(new_n654), .ZN(new_n748));
  OR3_X1    g562(.A1(new_n582), .A2(new_n294), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n667), .B1(new_n666), .B2(new_n657), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n665), .A2(new_n669), .A3(KEYINPUT104), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n747), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n582), .A2(new_n294), .A3(new_n748), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n668), .B2(new_n670), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n747), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n663), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n629), .A2(new_n566), .B1(new_n634), .B2(new_n295), .ZN(new_n759));
  AND4_X1   g573(.A1(KEYINPUT107), .A2(new_n626), .A3(new_n641), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n641), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n622), .B2(new_n625), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT107), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n530), .A2(new_n532), .ZN(new_n765));
  INV_X1    g579(.A(new_n436), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n577), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n229), .A2(new_n245), .B1(new_n547), .B2(new_n549), .ZN(new_n768));
  INV_X1    g582(.A(new_n294), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n612), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n256), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n435), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n560), .A3(new_n386), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT108), .ZN(new_n775));
  INV_X1    g589(.A(new_n773), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n533), .A2(new_n776), .A3(new_n577), .A4(KEYINPUT108), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n758), .A2(new_n764), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n746), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT53), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n746), .B2(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT112), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n741), .A2(new_n744), .A3(KEYINPUT52), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n626), .A2(new_n759), .A3(new_n641), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n762), .A2(KEYINPUT107), .A3(new_n759), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n767), .B2(new_n773), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n777), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n788), .A2(new_n797), .A3(new_n758), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n783), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n784), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n783), .B1(new_n656), .B2(new_n659), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n789), .B1(new_n753), .B2(new_n757), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n788), .A2(new_n779), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n798), .A2(KEYINPUT113), .A3(new_n783), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(new_n804), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n701), .A2(new_n536), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT115), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n716), .A2(new_n801), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(G952), .B2(G953), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n594), .A2(new_n673), .A3(new_n554), .A4(new_n297), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n620), .B(KEYINPUT49), .Z(new_n815));
  NAND4_X1  g629(.A1(new_n604), .A2(new_n434), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(G75));
  NAND3_X1  g631(.A1(new_n803), .A2(new_n807), .A3(new_n808), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(G210), .A3(G902), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n420), .A2(new_n425), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(new_n423), .Z(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT55), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n822), .A2(new_n825), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n189), .A2(G952), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G51));
  INV_X1    g643(.A(new_n663), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n756), .B1(new_n755), .B2(new_n747), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n791), .B(new_n792), .C1(new_n795), .C2(new_n777), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n802), .B(KEYINPUT53), .C1(new_n835), .C2(new_n788), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT113), .B1(new_n798), .B2(new_n783), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT117), .A3(new_n804), .A4(new_n807), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n809), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n379), .B(KEYINPUT57), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n382), .A2(new_n384), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n818), .A2(G469), .A3(G902), .A4(new_n678), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT118), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n828), .B1(new_n847), .B2(new_n849), .ZN(G54));
  AND3_X1   g664(.A1(new_n818), .A2(KEYINPUT58), .A3(G902), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(KEYINPUT119), .A3(G475), .A4(new_n242), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n818), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n854));
  INV_X1    g668(.A(new_n242), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n828), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n854), .A2(KEYINPUT120), .A3(new_n855), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT120), .B1(new_n854), .B2(new_n855), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n857), .A2(new_n861), .ZN(G60));
  XNOR2_X1  g676(.A(new_n548), .B(KEYINPUT59), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n801), .B2(new_n809), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n546), .B(KEYINPUT121), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n858), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n863), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n843), .B2(new_n868), .ZN(G63));
  NAND2_X1  g683(.A1(G217), .A2(G902), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT60), .Z(new_n871));
  NAND2_X1  g685(.A1(new_n818), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(new_n573), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n510), .A2(new_n511), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n858), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n873), .A2(KEYINPUT61), .A3(new_n858), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(G66));
  INV_X1    g694(.A(G224), .ZN(new_n881));
  OAI21_X1  g695(.A(G953), .B1(new_n254), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n797), .B2(G953), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n823), .B1(G898), .B2(new_n189), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(G69));
  XNOR2_X1  g699(.A(new_n463), .B(KEYINPUT122), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n235), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n685), .A2(new_n691), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n741), .B(new_n610), .C1(KEYINPUT123), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n606), .A2(new_n653), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n765), .A2(new_n770), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n741), .A2(new_n610), .ZN(new_n893));
  XOR2_X1   g707(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n888), .A2(new_n890), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n887), .B1(new_n896), .B2(new_n189), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n741), .A2(new_n671), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n684), .A2(new_n658), .A3(new_n722), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n888), .A2(new_n830), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n189), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n584), .B(KEYINPUT124), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n897), .B1(new_n904), .B2(new_n887), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n905), .B(new_n906), .Z(G72));
  XNOR2_X1  g721(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n557), .A2(new_n227), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT126), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n901), .B2(new_n834), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n466), .A2(new_n455), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n828), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT127), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n911), .B1(new_n896), .B2(new_n834), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n598), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n598), .A2(new_n913), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n785), .A2(new_n800), .A3(new_n910), .A4(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(G57));
endmodule


