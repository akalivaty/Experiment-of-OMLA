//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  OR2_X1    g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G43gat), .A2(G50gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  AOI211_X1 g012(.A(new_n204), .B(new_n208), .C1(new_n209), .C2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT94), .B(G43gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n205), .B(new_n207), .C1(new_n215), .C2(G50gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n216), .C1(new_n209), .C2(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n213), .A2(new_n218), .B1(new_n202), .B2(new_n203), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT93), .B1(new_n210), .B2(new_n212), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n223));
  XNOR2_X1  g022(.A(G99gat), .B(G106gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT104), .ZN(new_n225));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT7), .ZN(new_n227));
  INV_X1    g026(.A(G99gat), .ZN(new_n228));
  INV_X1    g027(.A(G106gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT8), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(new_n230), .C1(G85gat), .C2(G92gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n225), .B(new_n231), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n221), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT105), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n235), .A3(KEYINPUT105), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n233), .A2(new_n232), .B1(KEYINPUT41), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G190gat), .B(G218gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n240), .A2(new_n247), .A3(new_n243), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT106), .B1(new_n244), .B2(new_n245), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n242), .A2(KEYINPUT41), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G162gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n249), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n246), .A2(KEYINPUT106), .A3(new_n248), .A4(new_n254), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G71gat), .A2(G78gat), .ZN(new_n259));
  OR2_X1    g058(.A1(G71gat), .A2(G78gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G57gat), .B(G64gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT98), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT100), .ZN(new_n266));
  INV_X1    g065(.A(G57gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(G64gat), .ZN(new_n268));
  INV_X1    g067(.A(G64gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT99), .B(G57gat), .Z(new_n271));
  OAI211_X1 g070(.A(new_n268), .B(new_n270), .C1(new_n271), .C2(new_n269), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n260), .A2(new_n259), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT101), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n273), .A2(new_n274), .B1(new_n262), .B2(new_n259), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n275), .C1(new_n274), .C2(new_n273), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n265), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G127gat), .ZN(new_n282));
  XOR2_X1   g081(.A(G183gat), .B(G211gat), .Z(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G15gat), .B(G22gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT16), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(G1gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n289), .B(new_n290), .C1(G1gat), .C2(new_n287), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n277), .B2(new_n278), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(KEYINPUT103), .Z(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT102), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(G155gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n295), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n299), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n258), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n277), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n232), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n225), .B(new_n231), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n277), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n310), .B(KEYINPUT108), .Z(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(KEYINPUT107), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(KEYINPUT107), .A3(KEYINPUT10), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(new_n305), .A3(new_n309), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n311), .A2(new_n320), .A3(new_n316), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT97), .ZN(new_n327));
  XNOR2_X1  g126(.A(G15gat), .B(G43gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G71gat), .B(G99gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT66), .ZN(new_n332));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT24), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  OR3_X1    g137(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G169gat), .ZN(new_n341));
  INV_X1    g140(.A(G176gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT23), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(G169gat), .B2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT25), .A4(new_n346), .ZN(new_n349));
  INV_X1    g148(.A(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n337), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n332), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n352), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n347), .A3(KEYINPUT25), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n357));
  INV_X1    g156(.A(new_n338), .ZN(new_n358));
  NOR3_X1   g157(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n360), .B2(new_n337), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n356), .B(KEYINPUT66), .C1(new_n361), .C2(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  INV_X1    g164(.A(G120gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT73), .ZN(new_n367));
  OAI21_X1  g166(.A(G113gat), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT74), .B(KEYINPUT1), .Z(new_n369));
  INV_X1    g168(.A(G127gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G134gat), .ZN(new_n371));
  INV_X1    g170(.A(G113gat), .ZN(new_n372));
  INV_X1    g171(.A(G134gat), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n372), .A2(new_n366), .B1(new_n373), .B2(G127gat), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n368), .A2(new_n369), .A3(new_n371), .A4(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT1), .B1(new_n372), .B2(new_n366), .ZN(new_n376));
  NAND2_X1  g175(.A1(G113gat), .A2(G120gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(new_n373), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n370), .B2(G134gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n373), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n378), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n333), .ZN(new_n388));
  NOR2_X1   g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n346), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT69), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT26), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n395), .B2(KEYINPUT70), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT70), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n388), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n350), .A2(KEYINPUT27), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G183gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT68), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT27), .B(G183gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n351), .A2(KEYINPUT28), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n400), .A2(new_n402), .A3(new_n410), .A4(new_n351), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT28), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n406), .B2(new_n351), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n408), .A2(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n363), .A2(new_n387), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n387), .B1(new_n363), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n419), .B(KEYINPUT64), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n331), .B1(new_n422), .B2(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n363), .A2(new_n416), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n375), .A2(new_n386), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n354), .A2(new_n362), .B1(new_n415), .B2(new_n399), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n387), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n428), .A3(new_n420), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT75), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n331), .A2(KEYINPUT33), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(KEYINPUT32), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT76), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT76), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n429), .A2(new_n435), .A3(KEYINPUT32), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n330), .B1(new_n429), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n431), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT77), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n426), .A2(new_n446), .A3(new_n428), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n447), .A3(new_n419), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n420), .A2(KEYINPUT34), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n448), .A2(KEYINPUT34), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n450), .A2(new_n437), .A3(new_n431), .A4(new_n442), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT36), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n452), .A2(KEYINPUT78), .A3(KEYINPUT36), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n459), .A3(new_n453), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n443), .A2(KEYINPUT79), .A3(new_n451), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G57gat), .B(G85gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G225gat), .A2(G233gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G155gat), .A2(G162gat), .ZN(new_n471));
  INV_X1    g270(.A(G155gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n253), .ZN(new_n473));
  XNOR2_X1  g272(.A(G141gat), .B(G148gat), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n471), .B(new_n473), .C1(new_n474), .C2(KEYINPUT2), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n472), .A3(new_n253), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n471), .ZN(new_n478));
  INV_X1    g277(.A(G141gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(G148gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G148gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G141gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(G148gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT84), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n475), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n387), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n477), .A2(new_n471), .B1(new_n480), .B2(KEYINPUT84), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n386), .A2(new_n375), .B1(new_n493), .B2(new_n475), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n470), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT5), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT4), .B1(new_n387), .B2(new_n488), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n476), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n473), .A2(new_n471), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n492), .A2(new_n490), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n386), .A4(new_n375), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n425), .A2(new_n505), .A3(new_n502), .A4(new_n501), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(KEYINPUT4), .C1(new_n387), .C2(new_n488), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n498), .A2(new_n504), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n488), .A2(KEYINPUT3), .B1(new_n386), .B2(new_n375), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n470), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n496), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n503), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n468), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n513), .ZN(new_n519));
  INV_X1    g318(.A(new_n496), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  INV_X1    g321(.A(new_n468), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT89), .B(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n514), .A2(new_n468), .A3(new_n517), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n518), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n518), .A2(new_n526), .B1(new_n528), .B2(new_n525), .ZN(new_n529));
  XNOR2_X1  g328(.A(G197gat), .B(G204gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT22), .ZN(new_n531));
  INV_X1    g330(.A(G211gat), .ZN(new_n532));
  INV_X1    g331(.A(G218gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G211gat), .B(G218gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n539));
  NAND2_X1  g338(.A1(G226gat), .A2(G233gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n424), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT82), .B1(new_n427), .B2(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n340), .A2(new_n347), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n356), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n416), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n542), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n541), .A2(KEYINPUT29), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n424), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n416), .A2(new_n541), .A3(new_n547), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n535), .B(new_n536), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT80), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n553), .A2(KEYINPUT81), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n552), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n554), .B(new_n556), .C1(new_n427), .C2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT81), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n538), .A2(new_n551), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G8gat), .B(G36gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(G64gat), .B(G92gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(KEYINPUT30), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n538), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n557), .A2(new_n561), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT90), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n567), .A2(new_n568), .A3(new_n565), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n529), .A2(new_n572), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n521), .A2(new_n523), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n525), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR4_X1   g379(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n517), .A4(new_n468), .ZN(new_n581));
  INV_X1    g380(.A(new_n525), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n518), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n576), .A2(new_n566), .A3(new_n571), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT90), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G228gat), .ZN(new_n588));
  INV_X1    g387(.A(G233gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n512), .A2(new_n549), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n556), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n538), .A2(new_n549), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n501), .B1(new_n594), .B2(new_n511), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n555), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT31), .B(G50gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n600), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n604), .B2(new_n597), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G78gat), .B(G106gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G22gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n608), .A3(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n458), .A2(new_n463), .B1(new_n587), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n574), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n580), .B2(new_n583), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n565), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n569), .B2(new_n570), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n562), .A2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT38), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n542), .B(new_n555), .C1(new_n543), .C2(new_n550), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT91), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n399), .A2(new_n415), .B1(new_n546), .B2(new_n356), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n540), .B1(new_n623), .B2(KEYINPUT29), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n624), .B(KEYINPUT82), .C1(new_n540), .C2(new_n427), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n555), .A4(new_n542), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n553), .A2(new_n554), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n538), .B(KEYINPUT80), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n622), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT37), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n565), .B1(new_n562), .B2(new_n616), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n615), .A2(new_n620), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n510), .A2(new_n512), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n469), .B1(new_n516), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n468), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n387), .B(new_n488), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT39), .B1(new_n641), .B2(new_n470), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n645), .A2(new_n646), .A3(new_n579), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n612), .B1(new_n585), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n636), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT92), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n612), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n452), .A2(new_n654), .A3(new_n453), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT35), .B1(new_n587), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n460), .A2(new_n462), .ZN(new_n657));
  INV_X1    g456(.A(new_n585), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n657), .A2(new_n529), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n613), .A2(new_n653), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n233), .A2(new_n234), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n223), .A2(new_n293), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G229gat), .A2(G233gat), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n222), .A2(new_n293), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n663), .A2(KEYINPUT18), .A3(new_n664), .A4(new_n665), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n222), .B(new_n293), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n664), .B(KEYINPUT13), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G113gat), .B(G141gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G197gat), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT11), .B(G169gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT12), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n668), .A2(new_n680), .A3(new_n669), .A4(new_n672), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n327), .B1(new_n661), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n458), .A2(new_n463), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n577), .A2(new_n586), .A3(new_n612), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n653), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n656), .A2(new_n660), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(KEYINPUT97), .A3(new_n682), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n326), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n584), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  AND3_X1   g493(.A1(new_n691), .A2(new_n585), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G8gat), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n691), .B2(new_n585), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n691), .A2(new_n585), .A3(new_n694), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(G1325gat));
  AOI21_X1  g501(.A(G15gat), .B1(new_n691), .B2(new_n657), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n685), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n458), .A2(KEYINPUT109), .A3(new_n463), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G15gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT110), .Z(new_n709));
  AOI21_X1  g508(.A(new_n703), .B1(new_n691), .B2(new_n709), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n612), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NAND3_X1  g512(.A1(new_n258), .A2(new_n303), .A3(new_n325), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n684), .B2(new_n690), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n529), .A2(G29gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n303), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n683), .A3(new_n324), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n722));
  NAND2_X1  g521(.A1(new_n258), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n686), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n577), .A2(new_n586), .A3(KEYINPUT111), .A4(new_n612), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n705), .A2(new_n653), .A3(new_n706), .A4(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n723), .B1(new_n728), .B2(new_n688), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n689), .B2(new_n258), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n721), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G29gat), .B1(new_n732), .B2(new_n529), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n716), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n733), .A3(new_n734), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n715), .A2(new_n203), .A3(new_n585), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n732), .B2(new_n658), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n707), .A2(new_n215), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n721), .B(new_n742), .C1(new_n729), .C2(new_n731), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n715), .A2(new_n657), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n741), .B(new_n743), .C1(new_n744), .C2(new_n215), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n215), .B1(new_n715), .B2(new_n657), .ZN(new_n746));
  INV_X1    g545(.A(new_n743), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n612), .A2(G50gat), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n721), .B(new_n751), .C1(new_n729), .C2(new_n731), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n715), .A2(new_n612), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n750), .B(new_n752), .C1(new_n753), .C2(G50gat), .ZN(new_n754));
  AOI21_X1  g553(.A(G50gat), .B1(new_n715), .B2(new_n612), .ZN(new_n755));
  INV_X1    g554(.A(new_n752), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT48), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1331gat));
  NAND2_X1  g557(.A1(new_n728), .A2(new_n688), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n258), .A2(new_n303), .A3(new_n682), .A4(new_n325), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n584), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(new_n271), .ZN(G1332gat));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n585), .A3(new_n760), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT49), .B(G64gat), .Z(new_n766));
  OR2_X1    g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(new_n657), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n761), .A2(G71gat), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n707), .ZN(new_n776));
  OAI21_X1  g575(.A(G71gat), .B1(new_n761), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n775), .B2(new_n777), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n612), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n303), .A2(new_n683), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n303), .A2(KEYINPUT115), .A3(new_n683), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n258), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n759), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n792), .B(new_n789), .C1(new_n728), .C2(new_n688), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(G85gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n584), .A4(new_n324), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n729), .A2(new_n731), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n788), .B2(new_n324), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT116), .B(new_n325), .C1(new_n786), .C2(new_n787), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n584), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n796), .B1(new_n805), .B2(new_n795), .ZN(G1336gat));
  OAI211_X1 g605(.A(new_n585), .B(new_n801), .C1(new_n729), .C2(new_n731), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n325), .A2(G92gat), .A3(new_n658), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n791), .B2(new_n793), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1337gat));
  NAND4_X1  g614(.A1(new_n794), .A2(new_n228), .A3(new_n657), .A4(new_n324), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n803), .A2(new_n707), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n818), .B2(new_n228), .ZN(G1338gat));
  OAI211_X1 g618(.A(new_n612), .B(new_n801), .C1(new_n729), .C2(new_n731), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n324), .A2(new_n229), .A3(new_n612), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT117), .Z(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n791), .B2(new_n793), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1339gat));
  NAND3_X1  g628(.A1(new_n304), .A2(new_n683), .A3(new_n325), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n256), .A2(new_n257), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n670), .A2(new_n671), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n664), .B1(new_n663), .B2(new_n665), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n677), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n681), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n324), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  INV_X1    g636(.A(new_n305), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n315), .A2(new_n309), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT10), .B1(new_n307), .B2(KEYINPUT107), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n841), .A2(KEYINPUT54), .A3(new_n316), .ZN(new_n842));
  XOR2_X1   g641(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n321), .B1(new_n316), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n837), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(KEYINPUT54), .A3(new_n316), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n839), .A2(new_n840), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n305), .A3(new_n843), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT55), .A4(new_n321), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n323), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n836), .B1(new_n851), .B2(new_n683), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n256), .A2(new_n835), .A3(new_n257), .ZN(new_n853));
  INV_X1    g652(.A(new_n851), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n831), .A2(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n830), .B1(new_n855), .B2(new_n720), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n584), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(new_n585), .A3(new_n655), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n682), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n852), .A2(new_n831), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n854), .A2(new_n257), .A3(new_n256), .A4(new_n835), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n720), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n258), .A2(new_n303), .A3(new_n682), .A4(new_n324), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n657), .A2(new_n654), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n529), .A2(new_n585), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n372), .A3(new_n683), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n859), .A2(new_n869), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n868), .B2(new_n325), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n365), .A2(new_n367), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n858), .A2(new_n872), .A3(new_n324), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1341gat));
  OAI22_X1  g673(.A1(new_n868), .A2(new_n303), .B1(new_n380), .B2(new_n379), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n303), .A2(new_n380), .A3(new_n379), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1342gat));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n373), .A3(new_n258), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n868), .B2(new_n831), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  NOR3_X1   g682(.A1(new_n857), .A2(new_n585), .A3(new_n654), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n479), .A3(new_n682), .A4(new_n776), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n850), .A2(new_n323), .ZN(new_n887));
  INV_X1    g686(.A(new_n845), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT55), .B1(new_n888), .B2(new_n847), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n886), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n846), .A2(KEYINPUT119), .A3(new_n323), .A4(new_n850), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n682), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n258), .B1(new_n892), .B2(new_n836), .ZN(new_n893));
  INV_X1    g692(.A(new_n861), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n303), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n654), .B1(new_n895), .B2(new_n830), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n856), .A2(new_n897), .A3(new_n612), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n705), .A2(new_n706), .A3(new_n867), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n898), .A2(new_n901), .A3(new_n683), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n885), .B1(new_n902), .B2(new_n479), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(new_n885), .C1(new_n902), .C2(new_n479), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT57), .B(new_n612), .C1(new_n862), .C2(new_n863), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n856), .A2(new_n911), .A3(KEYINPUT57), .A4(new_n612), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n910), .B(new_n912), .C1(new_n896), .C2(KEYINPUT57), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n324), .A3(new_n900), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n908), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n901), .A3(new_n325), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(KEYINPUT59), .A3(new_n483), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n884), .A2(new_n776), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n324), .A2(new_n483), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n915), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1345gat));
  NOR4_X1   g719(.A1(new_n898), .A2(new_n901), .A3(new_n472), .A4(new_n303), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n918), .A2(new_n303), .ZN(new_n922));
  AOI21_X1  g721(.A(G155gat), .B1(new_n922), .B2(KEYINPUT121), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n918), .B2(new_n303), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n923), .B2(new_n925), .ZN(G1346gat));
  NAND4_X1  g725(.A1(new_n884), .A2(new_n253), .A3(new_n258), .A4(new_n776), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n898), .A2(new_n901), .A3(new_n831), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n253), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g730(.A(KEYINPUT122), .B(new_n927), .C1(new_n928), .C2(new_n253), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n658), .A2(new_n584), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n864), .A2(new_n865), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n683), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n935), .A2(new_n655), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n864), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n341), .A3(new_n682), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(G1348gat));
  NAND3_X1  g743(.A1(new_n936), .A2(G176gat), .A3(new_n324), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  AOI21_X1  g747(.A(G176gat), .B1(new_n940), .B2(new_n324), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n937), .B2(new_n303), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n303), .A2(new_n408), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT60), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n951), .B(new_n958), .C1(new_n954), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n940), .A2(new_n351), .A3(new_n258), .ZN(new_n961));
  OAI21_X1  g760(.A(G190gat), .B1(new_n937), .B2(new_n831), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1351gat));
  NOR2_X1   g764(.A1(new_n707), .A2(new_n935), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n913), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(G197gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n967), .A2(new_n968), .A3(new_n683), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n612), .A3(new_n856), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n970), .A2(new_n683), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(G1352gat));
  NAND3_X1  g771(.A1(new_n913), .A2(new_n324), .A3(new_n966), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G204gat), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n325), .A2(G204gat), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT62), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n970), .A2(KEYINPUT62), .A3(new_n975), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n974), .B(new_n976), .C1(new_n978), .C2(new_n979), .ZN(G1353gat));
  NAND3_X1  g779(.A1(new_n913), .A2(new_n720), .A3(new_n966), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G211gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT63), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n984), .A3(G211gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n720), .A2(new_n532), .ZN(new_n986));
  OR3_X1    g785(.A1(new_n970), .A2(KEYINPUT127), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT127), .B1(new_n970), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n983), .A2(new_n985), .A3(new_n989), .ZN(G1354gat));
  OAI21_X1  g789(.A(G218gat), .B1(new_n967), .B2(new_n831), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n258), .A2(new_n533), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n970), .B2(new_n992), .ZN(G1355gat));
endmodule


