//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n209));
  OR2_X1    g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT81), .ZN(new_n214));
  AND2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT79), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n221));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n217), .A2(new_n223), .A3(new_n212), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n211), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT80), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n214), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n208), .A2(KEYINPUT79), .B1(new_n211), .B2(new_n210), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n211), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(KEYINPUT81), .A3(new_n234), .A4(new_n223), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n213), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT22), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT72), .B(G211gat), .ZN(new_n238));
  INV_X1    g037(.A(G218gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G197gat), .B(G204gat), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n240), .A2(new_n242), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n244), .ZN(new_n248));
  INV_X1    g047(.A(G211gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT72), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G211gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT22), .B1(new_n253), .B2(G218gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n248), .B1(new_n254), .B2(new_n241), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n244), .A3(new_n242), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT85), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n236), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n228), .A2(new_n235), .ZN(new_n262));
  INV_X1    g061(.A(new_n213), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n264), .B2(new_n246), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n207), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT86), .B(new_n207), .C1(new_n260), .C2(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n207), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT29), .B1(new_n236), .B2(new_n259), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n255), .A2(KEYINPUT73), .A3(new_n256), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n236), .A2(new_n278), .ZN(new_n279));
  AOI211_X1 g078(.A(KEYINPUT82), .B(new_n213), .C1(new_n228), .C2(new_n235), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT3), .B1(new_n261), .B2(new_n246), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n206), .B1(new_n270), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g084(.A(G22gat), .B(new_n283), .C1(new_n268), .C2(new_n269), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n205), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n269), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT3), .B1(new_n247), .B2(new_n257), .ZN(new_n289));
  OAI22_X1  g088(.A1(new_n272), .A2(new_n261), .B1(new_n289), .B2(new_n236), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT86), .B1(new_n290), .B2(new_n207), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n284), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G22gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n270), .A2(new_n206), .A3(new_n284), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n204), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n276), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT27), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(G190gat), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT66), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n314), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(new_n312), .B2(new_n311), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n316), .A2(new_n319), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  INV_X1    g121(.A(G183gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n302), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n326), .A2(new_n331), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n336), .A2(new_n317), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(KEYINPUT25), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  INV_X1    g140(.A(new_n332), .ZN(new_n342));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n342), .A2(new_n333), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n336), .A2(new_n317), .A3(new_n338), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n321), .A2(new_n347), .A3(KEYINPUT74), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT74), .B1(new_n321), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n300), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n301), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n324), .B2(new_n325), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n302), .B1(new_n354), .B2(new_n307), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n316), .A2(new_n319), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n327), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n336), .A2(KEYINPUT25), .A3(new_n338), .A4(new_n317), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n304), .A2(new_n305), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n342), .B1(new_n361), .B2(new_n302), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n333), .B(new_n330), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n329), .B(new_n332), .C1(G183gat), .C2(G190gat), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT25), .B1(new_n339), .B2(new_n365), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n357), .A2(new_n359), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n299), .B1(new_n368), .B2(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n298), .B1(new_n351), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n348), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT75), .B1(new_n373), .B2(new_n300), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n297), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n246), .B1(new_n349), .B2(new_n350), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT76), .A3(new_n299), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n372), .B2(new_n348), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(new_n300), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n367), .A2(new_n300), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT77), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n377), .A2(new_n380), .A3(new_n261), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G8gat), .B(G36gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT78), .ZN(new_n386));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n383), .A3(new_n388), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT30), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n375), .A2(new_n383), .A3(new_n393), .A4(new_n388), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT40), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT67), .ZN(new_n398));
  INV_X1    g197(.A(G113gat), .ZN(new_n399));
  INV_X1    g198(.A(G120gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(G113gat), .B2(G120gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n398), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G127gat), .B(G134gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n264), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n236), .B(new_n278), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n259), .ZN(new_n410));
  INV_X1    g209(.A(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n236), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n236), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n397), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT39), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n412), .B1(new_n409), .B2(new_n411), .ZN(new_n427));
  INV_X1    g226(.A(new_n397), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT39), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n417), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n396), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n279), .A2(new_n280), .A3(new_n259), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n397), .B(new_n416), .C1(new_n432), .C2(new_n407), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n279), .A2(new_n280), .A3(new_n411), .ZN(new_n434));
  INV_X1    g233(.A(new_n412), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(KEYINPUT5), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT5), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n410), .A2(new_n438), .A3(new_n397), .A4(new_n416), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n424), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n424), .B1(new_n417), .B2(new_n418), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n442), .B(KEYINPUT40), .C1(new_n417), .C2(new_n429), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n431), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n296), .B1(new_n395), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n391), .ZN(new_n446));
  INV_X1    g245(.A(new_n374), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n351), .A2(new_n369), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n276), .C1(new_n448), .C2(new_n298), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n377), .A2(new_n380), .A3(new_n382), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(new_n261), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT38), .B1(new_n451), .B2(KEYINPUT37), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n389), .A2(KEYINPUT37), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n390), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n446), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n425), .A3(new_n439), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AND4_X1   g257(.A1(KEYINPUT84), .A2(new_n440), .A3(KEYINPUT6), .A4(new_n424), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n425), .B1(new_n437), .B2(new_n439), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT84), .B1(new_n460), .B2(KEYINPUT6), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n384), .A2(KEYINPUT37), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n389), .B1(new_n384), .B2(KEYINPUT37), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT38), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n455), .A2(new_n458), .A3(new_n462), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT87), .B1(new_n287), .B2(new_n295), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n295), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n441), .B2(new_n456), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n460), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n458), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n392), .A2(new_n394), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT70), .ZN(new_n479));
  NAND2_X1  g278(.A1(G227gat), .A2(G233gat), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n321), .A2(new_n347), .A3(new_n406), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n406), .B1(new_n321), .B2(new_n347), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT34), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n367), .A2(new_n411), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n321), .A2(new_n347), .A3(new_n406), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n480), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n484), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n484), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT68), .B(G71gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G99gat), .ZN(new_n495));
  XOR2_X1   g294(.A(G15gat), .B(G43gat), .Z(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n480), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n486), .A2(new_n498), .A3(new_n487), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(KEYINPUT32), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n499), .B(KEYINPUT32), .C1(new_n500), .C2(new_n497), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n479), .B1(new_n493), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n483), .A2(KEYINPUT34), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n489), .B1(new_n488), .B2(new_n480), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n503), .A3(new_n504), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT69), .B1(new_n508), .B2(new_n509), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n484), .A2(new_n485), .A3(new_n490), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n505), .A2(new_n479), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n507), .A2(KEYINPUT36), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n505), .B1(new_n509), .B2(new_n508), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n510), .A2(new_n503), .A3(new_n518), .A4(new_n504), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n467), .A2(new_n478), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n392), .B2(new_n394), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT35), .B1(new_n287), .B2(new_n295), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n526), .A2(new_n475), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n287), .A2(new_n295), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n511), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(new_n506), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n462), .A2(new_n458), .B1(new_n394), .B2(new_n392), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n531), .A3(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n528), .B1(new_n537), .B2(KEYINPUT35), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n525), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(G57gat), .A2(G64gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(G57gat), .A2(G64gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(KEYINPUT9), .ZN(new_n544));
  NOR2_X1   g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n542), .A2(new_n544), .B1(KEYINPUT95), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n543), .A2(new_n545), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT20), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n557), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n548), .A2(KEYINPUT98), .A3(new_n549), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT98), .B1(new_n548), .B2(new_n549), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT21), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G15gat), .B(G22gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(KEYINPUT91), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G1gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT16), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n571), .A3(new_n569), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(G8gat), .B1(new_n574), .B2(KEYINPUT92), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n573), .B(new_n574), .C1(KEYINPUT92), .C2(G8gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OR3_X1    g382(.A1(new_n562), .A2(new_n563), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n562), .B2(new_n563), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G36gat), .ZN(new_n590));
  AND2_X1   g389(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G29gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(KEYINPUT15), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(KEYINPUT15), .ZN(new_n598));
  XNOR2_X1  g397(.A(G43gat), .B(G50gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT17), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT17), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n577), .A2(KEYINPUT93), .A3(new_n578), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n577), .A2(new_n578), .A3(new_n602), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT18), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT90), .ZN(new_n616));
  XOR2_X1   g415(.A(G113gat), .B(G141gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G169gat), .B(G197gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n611), .A2(new_n612), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n610), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n602), .B1(new_n577), .B2(new_n578), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n609), .B(KEYINPUT13), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n614), .A2(new_n621), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n613), .A2(KEYINPUT18), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n621), .B1(new_n631), .B2(new_n623), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT101), .B(G85gat), .Z(new_n634));
  INV_X1    g433(.A(G92gat), .ZN(new_n635));
  INV_X1    g434(.A(G85gat), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT7), .B1(new_n636), .B2(new_n635), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT7), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(G85gat), .A3(G92gat), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n634), .A2(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT8), .ZN(new_n641));
  NAND2_X1  g440(.A1(G99gat), .A2(G106gat), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(KEYINPUT100), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(KEYINPUT100), .B2(new_n642), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G99gat), .B(G106gat), .Z(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT102), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n640), .A2(new_n647), .A3(new_n646), .A4(new_n644), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n606), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n653), .A2(new_n602), .B1(KEYINPUT41), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G190gat), .B(G218gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n662), .A3(new_n658), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n657), .A2(KEYINPUT41), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT99), .ZN(new_n665));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n661), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n661), .A2(KEYINPUT105), .A3(new_n663), .A4(new_n668), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT104), .B1(new_n659), .B2(new_n660), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n673), .A2(new_n663), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n667), .B1(new_n673), .B2(new_n663), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n671), .B(new_n672), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G230gat), .ZN(new_n677));
  INV_X1    g476(.A(G233gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n551), .A2(new_n653), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n645), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n646), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n645), .A2(new_n682), .A3(new_n649), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n550), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT10), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT10), .B(new_n653), .C1(new_n564), .C2(new_n565), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n680), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n550), .A2(new_n685), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n691), .A2(new_n684), .B1(new_n551), .B2(new_n653), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n679), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n690), .A2(new_n693), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR4_X1   g500(.A1(new_n587), .A2(new_n633), .A3(new_n676), .A4(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n539), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n475), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n462), .A2(KEYINPUT107), .A3(new_n458), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g509(.A1(new_n703), .A2(new_n395), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G8gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n711), .A2(KEYINPUT42), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT42), .B1(new_n711), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(G1325gat));
  INV_X1    g518(.A(new_n703), .ZN(new_n720));
  OAI21_X1  g519(.A(G15gat), .B1(new_n720), .B2(new_n524), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n520), .A2(G15gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(G1326gat));
  NAND2_X1  g522(.A1(new_n703), .A2(new_n471), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n676), .B1(new_n525), .B2(new_n538), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n633), .A2(new_n586), .A3(new_n701), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n708), .A2(new_n594), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n727), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n594), .A4(new_n708), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n523), .B1(new_n445), .B2(new_n466), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  INV_X1    g536(.A(new_n470), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n468), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n739), .B2(new_n535), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n471), .A2(KEYINPUT109), .A3(new_n477), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n743));
  INV_X1    g542(.A(new_n528), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT110), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n746), .B(new_n528), .C1(new_n537), .C2(KEYINPUT35), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n676), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(KEYINPUT44), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n748), .A2(new_n750), .B1(KEYINPUT44), .B2(new_n728), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n707), .A3(new_n730), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n734), .B(new_n735), .C1(new_n752), .C2(new_n594), .ZN(G1328gat));
  NAND2_X1  g552(.A1(new_n395), .A2(new_n590), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT46), .B1(new_n732), .B2(new_n754), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n751), .A2(new_n476), .A3(new_n730), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n590), .ZN(G1329gat));
  NAND2_X1  g557(.A1(new_n523), .A2(G43gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n751), .A2(new_n730), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n520), .ZN(new_n761));
  AOI21_X1  g560(.A(G43gat), .B1(new_n731), .B2(new_n761), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT47), .B1(new_n760), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1330gat));
  INV_X1    g564(.A(G50gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n471), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n732), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n748), .A2(new_n750), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n471), .B(new_n729), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n768), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n751), .A2(new_n730), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n766), .B1(new_n773), .B2(new_n296), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT48), .B1(new_n732), .B2(new_n767), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n772), .A2(KEYINPUT48), .B1(new_n774), .B2(new_n775), .ZN(G1331gat));
  AND3_X1   g575(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT35), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n529), .A2(KEYINPUT88), .A3(new_n531), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT88), .B1(new_n529), .B2(new_n531), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n778), .B1(new_n781), .B2(new_n535), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n746), .B1(new_n782), .B2(new_n528), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n538), .A2(KEYINPUT110), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n777), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n701), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n633), .A2(new_n586), .A3(new_n749), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n708), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g589(.A1(new_n476), .A2(new_n786), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n785), .A2(new_n787), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT49), .B(G64gat), .Z(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT111), .ZN(G1333gat));
  NAND2_X1  g598(.A1(new_n788), .A2(new_n523), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G71gat), .ZN(new_n801));
  INV_X1    g600(.A(G71gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n788), .A2(new_n802), .A3(new_n761), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n801), .A2(KEYINPUT50), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1334gat));
  NAND2_X1  g607(.A1(new_n788), .A2(new_n471), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G78gat), .ZN(G1335gat));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n587), .A2(new_n633), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n749), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n785), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n708), .A2(new_n634), .A3(new_n701), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n812), .A2(new_n786), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n751), .A2(new_n707), .A3(new_n821), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n818), .A2(new_n819), .B1(new_n822), .B2(new_n634), .ZN(G1336gat));
  NOR2_X1   g622(.A1(new_n792), .A2(G92gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n785), .A2(new_n811), .A3(new_n814), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n748), .B2(new_n813), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n751), .A2(new_n476), .A3(new_n821), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n635), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OAI221_X1 g632(.A(new_n827), .B1(new_n831), .B2(new_n830), .C1(new_n828), .C2(new_n635), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1337gat));
  INV_X1    g634(.A(G99gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n761), .A2(new_n836), .A3(new_n701), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n751), .A2(new_n524), .A3(new_n821), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n818), .A2(new_n837), .B1(new_n838), .B2(new_n836), .ZN(G1338gat));
  OAI211_X1 g638(.A(new_n471), .B(new_n820), .C1(new_n769), .C2(new_n770), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n529), .A2(G106gat), .A3(new_n786), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n840), .A2(G106gat), .B1(new_n817), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n817), .A2(new_n841), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n843), .ZN(new_n845));
  INV_X1    g644(.A(G106gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n751), .A2(new_n821), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n296), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n842), .A2(new_n843), .B1(new_n845), .B2(new_n848), .ZN(G1339gat));
  NAND4_X1  g648(.A1(new_n633), .A2(new_n586), .A3(new_n749), .A4(new_n786), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n679), .B(new_n688), .C1(new_n692), .C2(KEYINPUT10), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n690), .A2(new_n853), .A3(KEYINPUT54), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(new_n680), .C1(new_n687), .C2(new_n689), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n698), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n852), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n690), .A2(new_n853), .A3(KEYINPUT54), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(KEYINPUT55), .A3(new_n698), .A4(new_n856), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n700), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n621), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n614), .A2(new_n628), .ZN(new_n863));
  INV_X1    g662(.A(new_n623), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n865), .B2(new_n629), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n620), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT113), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n620), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n629), .A3(new_n701), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n749), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n858), .A2(new_n700), .A3(new_n860), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n676), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n629), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n851), .B1(new_n881), .B2(new_n587), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n707), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n476), .A3(new_n781), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n633), .ZN(new_n886));
  AOI21_X1  g685(.A(G113gat), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT114), .B1(new_n882), .B2(new_n471), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n877), .B1(new_n630), .B2(new_n632), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n676), .B1(new_n889), .B2(new_n874), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n878), .A2(new_n879), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n587), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n850), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n739), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n526), .A3(new_n708), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n633), .A2(new_n399), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n887), .B1(new_n898), .B2(new_n899), .ZN(G1340gat));
  AOI21_X1  g699(.A(G120gat), .B1(new_n885), .B2(new_n701), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n786), .A2(new_n400), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n898), .B2(new_n902), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n897), .B2(new_n587), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n587), .A2(G127gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n884), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n904), .B(KEYINPUT115), .C1(new_n884), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1342gat));
  NAND2_X1  g709(.A1(new_n883), .A2(new_n781), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n476), .A2(new_n676), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT116), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n911), .A2(G134gat), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g714(.A(G134gat), .B1(new_n897), .B2(new_n749), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1343gat));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n529), .B1(new_n892), .B2(new_n850), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT118), .B(new_n921), .C1(new_n882), .C2(new_n529), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n893), .A2(KEYINPUT57), .A3(new_n471), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n708), .A2(new_n476), .A3(new_n524), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT117), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G141gat), .B1(new_n927), .B2(new_n633), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n523), .A2(new_n529), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT119), .Z(new_n930));
  AND2_X1   g729(.A1(new_n883), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n476), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n218), .A3(new_n886), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT58), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n928), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1344gat));
  NAND2_X1  g737(.A1(new_n926), .A2(new_n701), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT57), .B1(new_n882), .B2(new_n529), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n893), .A2(new_n921), .A3(new_n471), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G148gat), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n701), .A3(new_n926), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n219), .A2(KEYINPUT59), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n219), .A3(new_n701), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1345gat));
  OAI21_X1  g751(.A(G155gat), .B1(new_n927), .B2(new_n587), .ZN(new_n953));
  INV_X1    g752(.A(G155gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n932), .A2(new_n954), .A3(new_n586), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1346gat));
  NOR2_X1   g755(.A1(new_n913), .A2(G162gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n931), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n959), .B1(new_n927), .B2(new_n749), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G162gat), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n927), .A2(new_n959), .A3(new_n749), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1347gat));
  AOI21_X1  g762(.A(new_n586), .B1(new_n876), .B2(new_n880), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n781), .B(new_n707), .C1(new_n964), .C2(new_n851), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n476), .ZN(new_n966));
  INV_X1    g765(.A(G169gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n886), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT122), .Z(new_n969));
  NAND3_X1  g768(.A1(new_n707), .A2(new_n395), .A3(new_n761), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n888), .B2(new_n895), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n967), .B1(new_n971), .B2(new_n886), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(G1348gat));
  INV_X1    g774(.A(new_n971), .ZN(new_n976));
  OAI21_X1  g775(.A(G176gat), .B1(new_n976), .B2(new_n786), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n792), .A2(G176gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n965), .B2(new_n978), .ZN(G1349gat));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980));
  INV_X1    g779(.A(new_n970), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n894), .B1(new_n893), .B2(new_n739), .ZN(new_n982));
  AOI211_X1 g781(.A(KEYINPUT114), .B(new_n471), .C1(new_n892), .C2(new_n850), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n586), .B(new_n981), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n361), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n586), .A2(new_n301), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n965), .A2(new_n476), .A3(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n980), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g789(.A(KEYINPUT125), .B(new_n988), .C1(new_n984), .C2(new_n985), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT60), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n992), .A2(KEYINPUT124), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n990), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n361), .B1(new_n971), .B2(new_n586), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n996), .B2(new_n988), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n986), .A2(new_n980), .A3(new_n989), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n995), .A2(new_n999), .ZN(G1350gat));
  NAND3_X1  g799(.A1(new_n966), .A2(new_n302), .A3(new_n676), .ZN(new_n1001));
  OAI21_X1  g800(.A(G190gat), .B1(new_n976), .B2(new_n749), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1002), .A2(KEYINPUT61), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1002), .A2(KEYINPUT61), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1351gat));
  NOR3_X1   g804(.A1(new_n708), .A2(new_n476), .A3(new_n523), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n940), .A2(new_n941), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(G197gat), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n1007), .A2(new_n1008), .A3(new_n633), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n882), .A2(new_n708), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1010), .A2(new_n395), .A3(new_n929), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n1011), .A2(new_n633), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1009), .B1(new_n1008), .B2(new_n1012), .ZN(G1352gat));
  NOR2_X1   g812(.A1(new_n792), .A2(G204gat), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1010), .A2(new_n929), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g814(.A(new_n1015), .B(KEYINPUT62), .Z(new_n1016));
  OAI21_X1  g815(.A(G204gat), .B1(new_n1007), .B2(new_n786), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1016), .A2(KEYINPUT126), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1020), .A2(new_n1021), .ZN(G1353gat));
  OR2_X1    g821(.A1(new_n1007), .A2(new_n587), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1023), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1023), .B2(G211gat), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n586), .A2(new_n238), .ZN(new_n1026));
  OAI22_X1  g825(.A1(new_n1024), .A2(new_n1025), .B1(new_n1011), .B2(new_n1026), .ZN(G1354gat));
  OAI21_X1  g826(.A(G218gat), .B1(new_n1007), .B2(new_n749), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n676), .A2(new_n239), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1028), .B1(new_n1011), .B2(new_n1029), .ZN(G1355gat));
endmodule


