//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G226gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n214), .C1(G169gat), .C2(G176gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT23), .B1(new_n216), .B2(KEYINPUT65), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n212), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n223));
  OR3_X1    g022(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n219), .B(KEYINPUT68), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n230), .A2(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n231), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n232), .A3(KEYINPUT25), .A4(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(KEYINPUT28), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n216), .B(KEYINPUT26), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n220), .B1(new_n239), .B2(new_n212), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n228), .A2(new_n234), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n209), .B1(new_n241), .B2(KEYINPUT29), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n228), .A2(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n208), .ZN(new_n246));
  XNOR2_X1  g045(.A(G197gat), .B(G204gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT22), .ZN(new_n248));
  INV_X1    g047(.A(G211gat), .ZN(new_n249));
  INV_X1    g048(.A(G218gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n242), .A2(new_n246), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n242), .B2(new_n246), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n205), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n208), .B1(new_n245), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n241), .A2(new_n209), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT30), .A3(new_n204), .A4(new_n256), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n204), .A3(new_n256), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT72), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G141gat), .B(G148gat), .Z(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT2), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G155gat), .B(G162gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n272), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n276), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT73), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n279), .A2(new_n272), .A3(KEYINPUT73), .A4(new_n275), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT3), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n285), .B2(new_n286), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n287), .C1(new_n285), .C2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n281), .A2(KEYINPUT3), .A3(new_n282), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n284), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n298));
  INV_X1    g097(.A(new_n293), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n292), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT69), .B1(new_n291), .B2(new_n292), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n298), .B(KEYINPUT4), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n295), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n281), .A2(new_n293), .A3(new_n282), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n309), .B2(new_n297), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n303), .A2(new_n304), .ZN(new_n312));
  INV_X1    g111(.A(new_n298), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n301), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n298), .A2(KEYINPUT4), .A3(new_n299), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n295), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT0), .ZN(new_n320));
  XNOR2_X1  g119(.A(G57gat), .B(G85gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n311), .A2(new_n322), .A3(new_n317), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n318), .A2(KEYINPUT6), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n271), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT81), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n259), .A2(new_n264), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n266), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n268), .ZN(new_n334));
  INV_X1    g133(.A(new_n329), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n254), .B1(new_n283), .B2(KEYINPUT29), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n254), .B2(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n313), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT74), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT76), .B(G22gat), .Z(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT75), .B(new_n254), .C1(new_n283), .C2(KEYINPUT29), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n340), .A4(new_n344), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n346), .A2(KEYINPUT77), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n354));
  AOI211_X1 g153(.A(new_n354), .B(new_n340), .C1(new_n341), .C2(new_n344), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n347), .B(new_n351), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n351), .B1(new_n353), .B2(new_n355), .ZN(new_n359));
  INV_X1    g158(.A(new_n347), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n352), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G78gat), .B(G106gat), .Z(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n356), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(G22gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n312), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n245), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n241), .A2(new_n312), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT34), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI211_X1 g177(.A(KEYINPUT34), .B(new_n372), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT70), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G71gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(G99gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n374), .A2(new_n372), .A3(new_n375), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(KEYINPUT32), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n385), .B(KEYINPUT32), .C1(new_n386), .C2(new_n384), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n380), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n378), .ZN(new_n393));
  INV_X1    g192(.A(new_n379), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n389), .A2(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT35), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n331), .A2(new_n338), .A3(new_n371), .A4(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT71), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT71), .B1(new_n378), .B2(new_n379), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n389), .A2(new_n390), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n392), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n336), .A2(new_n403), .A3(new_n371), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT35), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n366), .A2(new_n407), .A3(new_n370), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n366), .B2(new_n370), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n409), .A2(new_n410), .A3(new_n336), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n399), .A2(new_n400), .ZN(new_n412));
  INV_X1    g211(.A(new_n402), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT36), .B(new_n391), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT36), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n392), .B2(new_n395), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT37), .B1(new_n257), .B2(new_n258), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT37), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n263), .A2(new_n419), .A3(new_n256), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n205), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT79), .B(KEYINPUT38), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(KEYINPUT80), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(new_n205), .A3(new_n422), .A4(new_n420), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n426), .A2(new_n266), .A3(new_n327), .A4(new_n328), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT80), .B1(new_n421), .B2(new_n423), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT40), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n295), .A2(new_n314), .A3(new_n315), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n297), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n322), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n300), .A2(new_n296), .A3(new_n308), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT39), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n436), .B1(new_n431), .B2(new_n297), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n430), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n437), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT40), .A3(new_n322), .A4(new_n433), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n438), .A2(new_n440), .A3(new_n324), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n334), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n371), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n417), .B1(new_n429), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n406), .B1(new_n411), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G113gat), .B(G141gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT82), .B(G197gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT11), .B(G169gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT12), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  INV_X1    g252(.A(G43gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G50gat), .ZN(new_n455));
  INV_X1    g254(.A(G50gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G43gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT15), .ZN(new_n458));
  INV_X1    g257(.A(G29gat), .ZN(new_n459));
  INV_X1    g258(.A(G36gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT14), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(G29gat), .B2(G36gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n464), .A2(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n458), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n472), .A2(new_n458), .A3(new_n463), .A4(new_n461), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n454), .A2(KEYINPUT84), .A3(G50gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n453), .B1(new_n468), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT17), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n462), .A2(G29gat), .A3(G36gat), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT14), .B1(new_n459), .B2(new_n460), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT83), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G29gat), .A2(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n467), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n461), .A2(new_n491), .A3(new_n463), .A4(new_n469), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n488), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n477), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n475), .A3(new_n474), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(KEYINPUT86), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n481), .A2(new_n497), .A3(KEYINPUT87), .A4(new_n482), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(G1gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(new_n506), .C1(G1gat), .C2(new_n503), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n507), .B(G8gat), .Z(new_n508));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n487), .A2(new_n488), .B1(new_n493), .B2(new_n495), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(KEYINPUT17), .ZN(new_n511));
  AND4_X1   g310(.A1(new_n509), .A2(new_n489), .A3(KEYINPUT17), .A4(new_n496), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n502), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n508), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n481), .A2(new_n497), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n516), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n517), .B(new_n518), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n516), .B(KEYINPUT13), .Z(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n519), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n513), .B1(new_n500), .B2(new_n501), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(new_n508), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT18), .B1(new_n527), .B2(new_n516), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n452), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n520), .A3(new_n523), .A4(new_n451), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n445), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT41), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT94), .ZN(new_n539));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G85gat), .A2(G92gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT7), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  INV_X1    g349(.A(G92gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT96), .B1(new_n543), .B2(KEYINPUT7), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n543), .B2(new_n544), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n547), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT97), .ZN(new_n559));
  XOR2_X1   g358(.A(G99gat), .B(G106gat), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n553), .B2(new_n557), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n545), .A2(KEYINPUT7), .A3(new_n547), .ZN(new_n564));
  AND2_X1   g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n546), .B1(new_n565), .B2(new_n555), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(new_n561), .A3(new_n548), .A4(new_n552), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(KEYINPUT97), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n526), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G190gat), .B(G218gat), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n562), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n518), .A2(new_n573), .B1(KEYINPUT41), .B2(new_n537), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n570), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n542), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n571), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n541), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n584), .A2(KEYINPUT90), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n584), .B2(KEYINPUT90), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n583), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G64gat), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n592), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n593));
  INV_X1    g392(.A(G57gat), .ZN(new_n594));
  OR3_X1    g393(.A1(new_n594), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT91), .B1(new_n592), .B2(G57gat), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT92), .B1(new_n594), .B2(G64gat), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n593), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n583), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n589), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(G231gat), .B(G233gat), .C1(new_n602), .C2(KEYINPUT21), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G127gat), .ZN(new_n608));
  INV_X1    g407(.A(G127gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n517), .B1(KEYINPUT21), .B2(new_n602), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT93), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G155gat), .ZN(new_n618));
  XOR2_X1   g417(.A(G183gat), .B(G211gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n613), .A2(new_n614), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n569), .A2(new_n601), .A3(new_n562), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n563), .A2(new_n591), .A3(new_n600), .A4(new_n568), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n627), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n582), .A2(new_n624), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n535), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n335), .A2(KEYINPUT98), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n335), .A2(KEYINPUT98), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n334), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(G8gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G8gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT42), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(KEYINPUT42), .B2(new_n656), .ZN(G1325gat));
  INV_X1    g457(.A(new_n647), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n659), .B2(new_n417), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n392), .A2(new_n395), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(G15gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n660), .B1(new_n659), .B2(new_n663), .ZN(G1326gat));
  NOR2_X1   g463(.A1(new_n409), .A2(new_n410), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NOR3_X1   g467(.A1(new_n582), .A2(new_n624), .A3(new_n644), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n535), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n459), .A3(new_n650), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n396), .A2(new_n371), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n337), .B1(new_n271), .B2(new_n329), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n677), .A2(new_n338), .B1(KEYINPUT35), .B2(new_n404), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT101), .B1(new_n444), .B2(new_n411), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n334), .A2(new_n441), .B1(new_n366), .B2(new_n370), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n421), .A2(new_n423), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT80), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n327), .A2(new_n266), .A3(new_n328), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n683), .A2(new_n424), .A3(new_n426), .A4(new_n684), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n680), .A2(new_n685), .B1(new_n416), .B2(new_n414), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n330), .A3(new_n408), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n678), .B1(new_n679), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n674), .B1(new_n691), .B2(new_n582), .ZN(new_n692));
  INV_X1    g491(.A(new_n582), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n445), .A2(KEYINPUT44), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n624), .B(KEYINPUT99), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n644), .B(KEYINPUT100), .Z(new_n698));
  AND3_X1   g497(.A1(new_n697), .A2(new_n534), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n650), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n673), .A2(new_n702), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n670), .A2(G36gat), .A3(new_n271), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n700), .B2(new_n271), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(new_n454), .B1(new_n670), .B2(new_n662), .ZN(new_n708));
  INV_X1    g507(.A(new_n417), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n700), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1330gat));
  INV_X1    g512(.A(new_n371), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n692), .A2(new_n714), .A3(new_n694), .A4(new_n699), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n665), .A2(new_n456), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT103), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n671), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n719), .A3(KEYINPUT48), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n692), .A2(new_n665), .A3(new_n694), .A4(new_n699), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n719), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n720), .A2(new_n721), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n722), .A2(new_n727), .A3(new_n728), .ZN(G1331gat));
  NAND2_X1  g528(.A1(new_n680), .A2(new_n685), .ZN(new_n730));
  AND4_X1   g529(.A1(new_n687), .A2(new_n689), .A3(new_n730), .A4(new_n417), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n687), .B1(new_n686), .B2(new_n689), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n406), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n624), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n698), .A2(new_n693), .A3(new_n534), .A4(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n650), .B(KEYINPUT105), .Z(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g539(.A(new_n271), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  AOI21_X1  g547(.A(new_n587), .B1(new_n736), .B2(new_n709), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n662), .A2(G71gat), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n736), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n665), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n679), .A2(new_n690), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n582), .B1(new_n756), .B2(new_n406), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n534), .A2(new_n624), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT51), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  INV_X1    g559(.A(new_n758), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n691), .A2(new_n760), .A3(new_n582), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n755), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n733), .A2(new_n693), .A3(new_n758), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n760), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n693), .A4(new_n758), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(KEYINPUT110), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n701), .A2(G85gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n763), .A2(new_n644), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n758), .A2(new_n644), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT108), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n695), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n773), .B2(new_n701), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G85gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n770), .A3(new_n701), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  AOI21_X1  g576(.A(new_n698), .B1(new_n765), .B2(new_n766), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n551), .A3(new_n334), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n692), .A2(new_n334), .A3(new_n694), .A4(new_n772), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n779), .B(new_n781), .C1(new_n784), .C2(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1337gat));
  XNOR2_X1  g587(.A(KEYINPUT112), .B(G99gat), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n662), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n763), .A2(new_n644), .A3(new_n767), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n695), .A2(new_n709), .A3(new_n772), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n794), .A3(KEYINPUT113), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1338gat));
  OAI21_X1  g598(.A(G106gat), .B1(new_n773), .B2(new_n371), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n371), .A2(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n778), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n695), .A2(new_n665), .A3(new_n772), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n805), .A2(G106gat), .B1(new_n778), .B2(new_n801), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(G1339gat));
  NAND3_X1  g606(.A1(new_n582), .A2(new_n624), .A3(new_n645), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n534), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n516), .B1(new_n515), .B2(new_n519), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n521), .A2(new_n522), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n450), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT115), .B(new_n450), .C1(new_n810), .C2(new_n811), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n814), .A2(new_n533), .A3(new_n644), .A4(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n529), .A2(new_n533), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n640), .B1(new_n632), .B2(KEYINPUT54), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n628), .A2(new_n634), .A3(new_n629), .ZN(new_n821));
  AND4_X1   g620(.A1(new_n820), .A2(new_n632), .A3(KEYINPUT54), .A4(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n630), .B2(new_n631), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n820), .B1(new_n824), .B2(new_n821), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n819), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(KEYINPUT55), .B(new_n819), .C1(new_n822), .C2(new_n825), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n642), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n816), .B1(new_n817), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n830), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n533), .A3(new_n815), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n582), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n831), .A2(new_n582), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n696), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n824), .A2(new_n821), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n820), .A3(new_n821), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n818), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n641), .B1(new_n841), .B2(KEYINPUT55), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n534), .A2(new_n842), .A3(new_n828), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n693), .B1(new_n843), .B2(new_n816), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n830), .A2(new_n833), .A3(new_n582), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n809), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n737), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n403), .A2(new_n371), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(new_n271), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n534), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n847), .B2(new_n665), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n582), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n834), .A2(new_n832), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n836), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n846), .A3(new_n697), .ZN(new_n857));
  INV_X1    g656(.A(new_n809), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n665), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(KEYINPUT117), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n662), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n271), .A3(new_n650), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n817), .A2(new_n285), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n850), .B2(new_n644), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n698), .A2(new_n286), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n864), .B2(new_n868), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n863), .B2(new_n697), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n850), .A2(new_n609), .A3(new_n624), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n873), .A3(new_n693), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n863), .B2(new_n582), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NOR3_X1   g677(.A1(new_n701), .A2(new_n709), .A3(new_n334), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n371), .B1(new_n857), .B2(new_n858), .ZN(new_n880));
  XNOR2_X1  g679(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n665), .A2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n828), .A2(KEYINPUT119), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n826), .A2(new_n886), .A3(new_n827), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n534), .A2(new_n842), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n816), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n845), .B1(new_n890), .B2(new_n582), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(new_n624), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(new_n858), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n879), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894), .B2(new_n817), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n709), .A2(new_n334), .A3(new_n371), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n848), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n817), .A2(G141gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n895), .B(new_n901), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n646), .B2(new_n817), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n808), .A2(KEYINPUT122), .A3(new_n534), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n891), .B2(new_n624), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n665), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n880), .B2(new_n882), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n879), .A2(new_n644), .ZN(new_n912));
  OAI21_X1  g711(.A(G148gat), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n644), .B(new_n879), .C1(new_n883), .C2(new_n893), .ZN(new_n916));
  INV_X1    g715(.A(G148gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(KEYINPUT59), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n913), .A2(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n645), .A2(G148gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n848), .A2(new_n896), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n904), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n921), .B(KEYINPUT120), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n916), .A2(new_n918), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n847), .A2(new_n371), .A3(new_n881), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n644), .B(new_n879), .C1(new_n927), .C2(new_n910), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n914), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT123), .B(new_n925), .C1(new_n926), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n924), .A2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n894), .B2(new_n697), .ZN(new_n932));
  INV_X1    g731(.A(new_n897), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n273), .A3(new_n624), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n894), .B2(new_n582), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n274), .A3(new_n693), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1347gat));
  NOR3_X1   g737(.A1(new_n847), .A2(new_n271), .A3(new_n650), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n849), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n534), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n738), .A2(new_n271), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT117), .B1(new_n859), .B2(new_n860), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n852), .B(new_n665), .C1(new_n857), .C2(new_n858), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n661), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n534), .A2(G169gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(G1348gat));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950));
  INV_X1    g749(.A(G176gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n698), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n862), .A2(KEYINPUT124), .A3(new_n943), .A4(new_n952), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n940), .B2(new_n645), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n954), .A2(KEYINPUT125), .A3(new_n955), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1349gat));
  OAI21_X1  g760(.A(G183gat), .B1(new_n946), .B2(new_n697), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n941), .A2(new_n235), .A3(new_n624), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT60), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(KEYINPUT60), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n941), .A2(new_n236), .A3(new_n693), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n862), .A2(new_n693), .A3(new_n943), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(G190gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n971), .B2(G190gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  AND3_X1   g774(.A1(new_n939), .A2(new_n714), .A3(new_n417), .ZN(new_n976));
  XOR2_X1   g775(.A(KEYINPUT127), .B(G197gat), .Z(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(new_n534), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n943), .A2(new_n417), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n911), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n980), .A2(new_n817), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n981), .B2(new_n977), .ZN(G1352gat));
  INV_X1    g781(.A(G204gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n976), .A2(new_n983), .A3(new_n644), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n985));
  OAI21_X1  g784(.A(G204gat), .B1(new_n980), .B2(new_n698), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(G1353gat));
  NAND3_X1  g787(.A1(new_n976), .A2(new_n249), .A3(new_n624), .ZN(new_n989));
  OR3_X1    g788(.A1(new_n911), .A2(new_n734), .A3(new_n979), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  OAI21_X1  g792(.A(G218gat), .B1(new_n980), .B2(new_n582), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n250), .A3(new_n693), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


