//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(KEYINPUT75), .B2(KEYINPUT22), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT76), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT22), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(new_n213), .B1(G211gat), .B2(G218gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(new_n209), .ZN(new_n216));
  XNOR2_X1  g015(.A(G197gat), .B(G204gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G211gat), .B(G218gat), .Z(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n219), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n211), .A2(new_n221), .A3(new_n216), .A4(new_n217), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT79), .B(KEYINPUT2), .Z(new_n233));
  INV_X1    g032(.A(G162gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G155gat), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G162gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n232), .A2(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(KEYINPUT80), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G155gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(G162gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n235), .A3(new_n237), .A4(new_n231), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT80), .B(G155gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT2), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  AND4_X1   g049(.A1(new_n235), .A2(new_n230), .A3(new_n237), .A4(new_n231), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT81), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n239), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n227), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n224), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n226), .B(new_n239), .C1(new_n248), .C2(new_n252), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n246), .B1(new_n245), .B2(new_n247), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT81), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n238), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT82), .A3(new_n226), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n255), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n254), .B1(new_n263), .B2(new_n223), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n256), .A2(new_n257), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT82), .B1(new_n261), .B2(new_n226), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n224), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n220), .A2(new_n222), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n226), .B1(new_n268), .B2(KEYINPUT29), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n205), .B1(new_n270), .B2(new_n253), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n205), .A2(new_n264), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G22gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n271), .B1(new_n223), .B2(new_n263), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n261), .B1(new_n225), .B2(new_n226), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n267), .B2(new_n268), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n277), .B(new_n273), .C1(new_n279), .C2(new_n204), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(new_n275), .A3(new_n273), .ZN(new_n282));
  XNOR2_X1  g081(.A(G78gat), .B(G106gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT31), .B(G50gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  AND2_X1   g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT88), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT86), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n272), .B2(new_n273), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(KEYINPUT87), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT87), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n292), .A3(new_n273), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n285), .B1(new_n274), .B2(KEYINPUT86), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n277), .B1(new_n279), .B2(new_n204), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(KEYINPUT86), .A3(G22gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n285), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n297), .A2(new_n301), .A3(KEYINPUT88), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n287), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT34), .ZN(new_n304));
  INV_X1    g103(.A(G227gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(new_n203), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n310));
  INV_X1    g109(.A(G134gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(G127gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n309), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G113gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n311), .A2(G127gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n308), .A2(G134gat), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n323), .A2(new_n316), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n322), .A2(new_n326), .A3(KEYINPUT69), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT69), .B1(new_n322), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT70), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT70), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n326), .A3(KEYINPUT69), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G169gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n338), .A2(KEYINPUT26), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n339), .A2(KEYINPUT26), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G183gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G183gat), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G190gat), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT28), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n348), .A2(G183gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n346), .A2(KEYINPUT27), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT65), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G190gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n360), .B2(KEYINPUT66), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n356), .A2(new_n362), .A3(new_n357), .A4(new_n359), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n345), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT64), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT24), .B1(new_n341), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n365), .B2(new_n341), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n351), .ZN(new_n368));
  NAND3_X1  g167(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n336), .A2(new_n337), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n338), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n339), .A2(KEYINPUT23), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n373), .A2(KEYINPUT25), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n342), .A2(KEYINPUT24), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(new_n369), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n373), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n370), .A2(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n329), .B(new_n335), .C1(new_n364), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n360), .A2(KEYINPUT66), .ZN(new_n382));
  INV_X1    g181(.A(new_n352), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n363), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n344), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n332), .A2(new_n334), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n370), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n378), .A2(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n385), .A2(KEYINPUT70), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n306), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n304), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT73), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n390), .ZN(new_n397));
  INV_X1    g196(.A(new_n306), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n396), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n395), .B1(new_n391), .B2(new_n392), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n393), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT32), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n381), .A2(new_n390), .A3(new_n306), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n381), .A2(new_n390), .A3(KEYINPUT71), .A4(new_n306), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT33), .B1(new_n408), .B2(new_n409), .ZN(new_n411));
  XOR2_X1   g210(.A(G15gat), .B(G43gat), .Z(new_n412));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  AOI221_X4 g215(.A(new_n405), .B1(KEYINPUT33), .B2(new_n414), .C1(new_n408), .C2(new_n409), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n401), .B(new_n404), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n404), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n411), .A2(new_n415), .ZN(new_n420));
  INV_X1    g219(.A(new_n410), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n417), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n364), .B2(new_n380), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n385), .B2(new_n389), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT78), .B(new_n433), .C1(new_n434), .C2(new_n432), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n433), .A2(KEYINPUT78), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n268), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n364), .A2(new_n380), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n438), .B2(new_n255), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n223), .B1(new_n439), .B2(new_n433), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n430), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n433), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n268), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n433), .A2(KEYINPUT78), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n433), .A2(KEYINPUT78), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n431), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n443), .B(new_n429), .C1(new_n447), .C2(new_n268), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(new_n448), .A3(KEYINPUT30), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n437), .A2(new_n440), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n429), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT35), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT5), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n327), .A2(new_n328), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n261), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n258), .A2(new_n262), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n330), .B1(new_n261), .B2(new_n226), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT4), .B1(new_n386), .B2(new_n253), .ZN(new_n466));
  INV_X1    g265(.A(new_n330), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n261), .A2(new_n457), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(KEYINPUT84), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n461), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n463), .B1(new_n258), .B2(new_n262), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n457), .B1(new_n386), .B2(new_n253), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n467), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n456), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G225gat), .A2(G233gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT83), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n470), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n253), .A2(new_n330), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n261), .A2(new_n467), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT5), .A4(new_n477), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT90), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT0), .ZN(new_n486));
  XNOR2_X1  g285(.A(G57gat), .B(G85gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(KEYINPUT90), .A3(new_n482), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n479), .A2(new_n482), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n489), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AND4_X1   g295(.A1(KEYINPUT91), .A2(new_n493), .A3(KEYINPUT6), .A4(new_n489), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n488), .B1(new_n479), .B2(new_n482), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT91), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n455), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n303), .A2(new_n426), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT92), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n303), .A2(new_n501), .A3(new_n504), .A4(new_n426), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n418), .A2(new_n424), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n419), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(KEYINPUT74), .C1(new_n416), .C2(new_n417), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n303), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT93), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n494), .B2(new_n498), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n453), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n303), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n513), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n506), .B1(KEYINPUT35), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n516), .B(new_n287), .C1(new_n296), .C2(new_n302), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n449), .A2(new_n452), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT40), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT39), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n477), .C1(new_n471), .C2(new_n474), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n488), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n480), .A2(new_n481), .A3(new_n478), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT39), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT4), .B1(new_n458), .B2(new_n261), .ZN(new_n530));
  INV_X1    g329(.A(new_n473), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n465), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n533), .B2(new_n477), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n524), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT89), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(new_n524), .C1(new_n527), .C2(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n527), .A2(new_n534), .A3(new_n524), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n523), .A2(new_n491), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n514), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n498), .A2(KEYINPUT91), .A3(KEYINPUT6), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n479), .A2(KEYINPUT90), .A3(new_n482), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n545), .A2(new_n483), .A3(new_n488), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n543), .B(new_n544), .C1(new_n546), .C2(new_n494), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n429), .B1(new_n450), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n435), .A2(new_n436), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n268), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n442), .B2(new_n223), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT38), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n549), .A2(new_n553), .B1(new_n450), .B2(new_n429), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n443), .B1(new_n447), .B2(new_n268), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n430), .B1(new_n555), .B2(KEYINPUT37), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n450), .A2(new_n548), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT38), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n541), .B1(new_n547), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n291), .A2(new_n293), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(new_n295), .A3(new_n288), .A4(new_n290), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT88), .B1(new_n297), .B2(new_n301), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n562), .A2(new_n563), .B1(new_n281), .B2(new_n286), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n522), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT36), .B1(new_n418), .B2(new_n424), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n511), .B2(KEYINPUT36), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n521), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT94), .B(KEYINPUT12), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT95), .B(G36gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G29gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT14), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(KEYINPUT14), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT15), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n577), .A2(KEYINPUT15), .A3(new_n579), .A4(new_n580), .ZN(new_n584));
  XNOR2_X1  g383(.A(G43gat), .B(G50gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G15gat), .B(G22gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(G8gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT16), .ZN(new_n594));
  AOI21_X1  g393(.A(G1gat), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n589), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT13), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n598), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n589), .A2(new_n596), .ZN(new_n602));
  INV_X1    g401(.A(new_n596), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT17), .B1(new_n586), .B2(new_n587), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT97), .B1(new_n588), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n586), .A2(new_n587), .A3(new_n608), .A4(KEYINPUT17), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI211_X1 g409(.A(new_n601), .B(new_n602), .C1(new_n605), .C2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n600), .B1(new_n611), .B2(KEYINPUT18), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n602), .B1(new_n605), .B2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n598), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n575), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(KEYINPUT18), .ZN(new_n619));
  INV_X1    g418(.A(new_n575), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n600), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n569), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n626));
  XOR2_X1   g425(.A(G57gat), .B(G64gat), .Z(new_n627));
  INV_X1    g426(.A(KEYINPUT9), .ZN(new_n628));
  INV_X1    g427(.A(G71gat), .ZN(new_n629));
  INV_X1    g428(.A(G78gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G71gat), .B(G78gat), .Z(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n626), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n627), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n638));
  INV_X1    g437(.A(new_n633), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(KEYINPUT99), .A3(new_n634), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G127gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n596), .B1(new_n642), .B2(new_n643), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT100), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n647), .A2(new_n649), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n236), .ZN(new_n654));
  XOR2_X1   g453(.A(G183gat), .B(G211gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G85gat), .ZN(new_n660));
  INV_X1    g459(.A(G92gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n663));
  OR2_X1    g462(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G99gat), .A2(G106gat), .ZN(new_n666));
  AOI22_X1  g465(.A1(KEYINPUT8), .A2(new_n666), .B1(new_n660), .B2(new_n661), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n665), .B(new_n667), .C1(new_n662), .C2(new_n664), .ZN(new_n668));
  XOR2_X1   g467(.A(G99gat), .B(G106gat), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n668), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n604), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n610), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(G232gat), .A2(G233gat), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n588), .A2(new_n671), .B1(KEYINPUT41), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(G190gat), .B(G218gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n674), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(G134gat), .B(G162gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n678), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n625), .B1(new_n659), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n657), .A2(KEYINPUT102), .A3(new_n658), .A4(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n637), .A2(new_n671), .A3(KEYINPUT10), .A4(new_n641), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n668), .B(new_n669), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n637), .A2(new_n689), .A3(new_n641), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n640), .A2(new_n634), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT10), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT103), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n696), .B(KEYINPUT10), .C1(new_n690), .C2(new_n692), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n688), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(G230gat), .A2(G233gat), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n698), .A2(KEYINPUT104), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT104), .B1(new_n698), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n693), .A2(new_n699), .ZN(new_n703));
  XNOR2_X1  g502(.A(G120gat), .B(G148gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(G176gat), .B(G204gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n699), .B(KEYINPUT105), .Z(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n698), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n706), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n687), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n624), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n515), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g518(.A1(new_n624), .A2(new_n715), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n453), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n592), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT16), .B(G8gat), .Z(new_n723));
  AND3_X1   g522(.A1(new_n716), .A2(new_n523), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT42), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n723), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(G1325gat));
  OR3_X1    g528(.A1(new_n720), .A2(G15gat), .A3(new_n425), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n511), .A2(KEYINPUT36), .ZN(new_n731));
  INV_X1    g530(.A(new_n566), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G15gat), .B1(new_n720), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(G1326gat));
  XOR2_X1   g534(.A(KEYINPUT43), .B(G22gat), .Z(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n716), .A2(new_n564), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n720), .B2(new_n303), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(G1327gat));
  INV_X1    g542(.A(new_n659), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n714), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n684), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n624), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n515), .A2(G29gat), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n683), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n521), .B2(new_n568), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n617), .A2(KEYINPUT108), .A3(new_n621), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT108), .B1(new_n617), .B2(new_n621), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n744), .A2(new_n714), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n564), .A2(new_n425), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n504), .B1(new_n760), .B2(new_n501), .ZN(new_n761));
  INV_X1    g560(.A(new_n505), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n303), .A2(new_n511), .A3(new_n518), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n518), .B1(new_n303), .B2(new_n511), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n516), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n766), .B2(new_n454), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n565), .B2(new_n567), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n496), .A2(new_n500), .A3(new_n558), .A4(new_n554), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n303), .A2(new_n770), .A3(new_n541), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n733), .A2(KEYINPUT109), .A3(new_n771), .A4(new_n522), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n683), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n754), .B(new_n759), .C1(new_n774), .C2(KEYINPUT44), .ZN(new_n775));
  OAI21_X1  g574(.A(G29gat), .B1(new_n775), .B2(new_n515), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n751), .A2(new_n776), .A3(new_n777), .ZN(G1328gat));
  XNOR2_X1  g577(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n453), .A2(new_n576), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n748), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n576), .B1(new_n775), .B2(new_n453), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n748), .B2(new_n780), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(G1329gat));
  OAI21_X1  g583(.A(G43gat), .B1(new_n775), .B2(new_n733), .ZN(new_n785));
  INV_X1    g584(.A(G43gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n426), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g586(.A1(new_n569), .A2(new_n623), .A3(new_n746), .A4(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT47), .B1(new_n790), .B2(KEYINPUT111), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n772), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n684), .B1(new_n521), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n752), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n794), .A2(new_n567), .A3(new_n754), .A4(new_n759), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n788), .B1(new_n795), .B2(G43gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n791), .A2(new_n799), .ZN(G1330gat));
  INV_X1    g599(.A(G50gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n748), .B2(new_n303), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n564), .A2(G50gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n775), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT48), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT48), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n802), .B(new_n806), .C1(new_n775), .C2(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1331gat));
  NAND2_X1  g607(.A1(new_n758), .A2(new_n714), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n687), .B(new_n809), .C1(new_n767), .C2(new_n773), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n717), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g611(.A(new_n453), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(new_n816), .A3(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1333gat));
  NAND3_X1  g619(.A1(new_n810), .A2(new_n629), .A3(new_n426), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n810), .A2(new_n567), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n823), .B2(new_n629), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(G1334gat));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n564), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT113), .B(G78gat), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n827), .B(new_n828), .ZN(G1335gat));
  NOR2_X1   g628(.A1(new_n744), .A2(new_n809), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n794), .A2(new_n754), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G85gat), .B1(new_n831), .B2(new_n515), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n744), .A2(new_n757), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n774), .A2(KEYINPUT51), .A3(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n684), .B(new_n833), .C1(new_n521), .C2(new_n792), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n714), .A2(new_n660), .A3(new_n717), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT114), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n832), .B1(new_n838), .B2(new_n840), .ZN(G1336gat));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n837), .A3(KEYINPUT115), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n835), .A2(new_n843), .A3(new_n836), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n713), .A2(G92gat), .A3(new_n453), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G92gat), .B1(new_n831), .B2(new_n453), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n837), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(new_n850), .B2(new_n845), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n847), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(G1337gat));
  OAI21_X1  g652(.A(G99gat), .B1(new_n831), .B2(new_n733), .ZN(new_n854));
  OR3_X1    g653(.A1(new_n713), .A2(new_n425), .A3(G99gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n838), .B2(new_n855), .ZN(G1338gat));
  NOR3_X1   g655(.A1(new_n303), .A2(G106gat), .A3(new_n713), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n844), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G106gat), .B1(new_n831), .B2(new_n303), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT53), .B1(new_n850), .B2(new_n857), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1339gat));
  XOR2_X1   g663(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n865));
  NOR2_X1   g664(.A1(new_n711), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n706), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n700), .B2(new_n701), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n709), .B(new_n688), .C1(new_n695), .C2(new_n697), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT116), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n708), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n867), .B(KEYINPUT55), .C1(new_n868), .C2(new_n870), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n613), .A2(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n573), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n621), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n683), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n873), .A2(KEYINPUT118), .A3(new_n878), .A4(new_n874), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n873), .A2(new_n757), .A3(new_n874), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n713), .A2(new_n877), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n684), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n659), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n685), .A2(new_n686), .A3(new_n713), .A4(new_n758), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n515), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n764), .A2(new_n765), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n453), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n889), .A2(new_n453), .A3(new_n890), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n317), .A3(new_n757), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n887), .A2(new_n888), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n898), .A2(new_n717), .A3(new_n453), .A4(new_n760), .ZN(new_n899));
  OAI21_X1  g698(.A(G113gat), .B1(new_n899), .B2(new_n623), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(G1340gat));
  AOI211_X1 g700(.A(G120gat), .B(new_n713), .C1(new_n892), .C2(new_n895), .ZN(new_n902));
  INV_X1    g701(.A(new_n899), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n319), .B1(new_n903), .B2(new_n714), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n713), .A2(G120gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n896), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(G1341gat));
  OAI21_X1  g709(.A(G127gat), .B1(new_n899), .B2(new_n659), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n744), .A2(new_n308), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n893), .B2(new_n912), .ZN(G1342gat));
  NAND4_X1  g712(.A1(new_n891), .A2(new_n311), .A3(new_n453), .A4(new_n684), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g714(.A(G134gat), .B1(new_n899), .B2(new_n683), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G1343gat));
  NAND2_X1  g717(.A1(new_n871), .A2(new_n872), .ZN(new_n919));
  INV_X1    g718(.A(new_n708), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n622), .A3(new_n920), .A4(new_n874), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n684), .B1(new_n921), .B2(new_n885), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n659), .B1(new_n883), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n888), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT57), .B1(new_n924), .B2(new_n303), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n898), .A2(new_n926), .A3(new_n564), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n567), .A2(new_n515), .A3(new_n523), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n623), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(KEYINPUT58), .A3(new_n228), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n567), .A2(new_n303), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n889), .A2(new_n933), .ZN(new_n934));
  NOR4_X1   g733(.A1(new_n934), .A2(G141gat), .A3(new_n523), .A4(new_n623), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n925), .A2(new_n757), .A3(new_n927), .A4(new_n928), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n935), .A2(new_n939), .B1(new_n940), .B2(G141gat), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n931), .A2(new_n938), .B1(new_n941), .B2(new_n936), .ZN(G1344gat));
  NAND4_X1  g741(.A1(new_n925), .A2(new_n714), .A3(new_n927), .A4(new_n928), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n229), .A2(KEYINPUT59), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  INV_X1    g746(.A(new_n879), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n659), .B1(new_n922), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n685), .A2(new_n623), .A3(new_n686), .A4(new_n713), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n303), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n951), .A2(KEYINPUT124), .A3(KEYINPUT57), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n898), .A2(KEYINPUT57), .A3(new_n564), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT124), .B1(new_n951), .B2(KEYINPUT57), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n928), .A2(new_n714), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n229), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT59), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n946), .A2(new_n947), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n934), .A2(new_n523), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n229), .A3(new_n714), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1345gat));
  OAI21_X1  g762(.A(new_n244), .B1(new_n929), .B2(new_n659), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(new_n249), .A3(new_n744), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1346gat));
  OAI21_X1  g765(.A(G162gat), .B1(new_n929), .B2(new_n683), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n684), .A2(new_n234), .A3(new_n453), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n934), .B2(new_n968), .ZN(G1347gat));
  AOI21_X1  g768(.A(new_n717), .B1(new_n887), .B2(new_n888), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(new_n523), .A3(new_n890), .ZN(new_n971));
  AOI21_X1  g770(.A(G169gat), .B1(new_n971), .B2(new_n757), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n717), .A2(new_n453), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n898), .A2(new_n760), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n623), .A2(new_n336), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1348gat));
  INV_X1    g775(.A(new_n974), .ZN(new_n977));
  OAI21_X1  g776(.A(G176gat), .B1(new_n977), .B2(new_n713), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n971), .A2(new_n337), .A3(new_n714), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1349gat));
  AOI21_X1  g779(.A(new_n346), .B1(new_n974), .B2(new_n744), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n744), .A2(new_n356), .A3(new_n357), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n971), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n983), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g783(.A(new_n351), .B1(new_n974), .B2(new_n684), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT61), .Z(new_n986));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n351), .A3(new_n684), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1351gat));
  NAND2_X1  g787(.A1(new_n733), .A2(new_n973), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n954), .A2(new_n953), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n951), .A2(KEYINPUT124), .A3(KEYINPUT57), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n622), .B(new_n990), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(G197gat), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n970), .A2(new_n523), .A3(new_n932), .ZN(new_n995));
  INV_X1    g794(.A(G197gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n995), .A2(new_n996), .A3(new_n757), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n994), .A2(new_n1000), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n999), .A2(new_n1001), .ZN(G1352gat));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n955), .A2(new_n990), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n1004), .B2(new_n713), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n955), .A2(KEYINPUT127), .A3(new_n714), .A4(new_n990), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1005), .A2(G204gat), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(G204gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n995), .A2(new_n1008), .A3(new_n714), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  NAND2_X1  g809(.A1(new_n1007), .A2(new_n1010), .ZN(G1353gat));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n206), .A3(new_n744), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n991), .A2(new_n992), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n733), .A2(new_n744), .A3(new_n973), .ZN(new_n1014));
  OAI21_X1  g813(.A(G211gat), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT63), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1012), .B1(new_n1017), .B2(new_n1018), .ZN(G1354gat));
  NOR3_X1   g818(.A1(new_n1004), .A2(new_n207), .A3(new_n683), .ZN(new_n1020));
  AOI21_X1  g819(.A(G218gat), .B1(new_n995), .B2(new_n684), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n1020), .A2(new_n1021), .ZN(G1355gat));
endmodule


