//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G137), .A4(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n467), .B2(new_n468), .ZN(new_n476));
  AND2_X1   g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT69), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n469), .A2(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n483), .B(new_n486), .C1(G136), .C2(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT70), .B(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n496), .B(new_n500), .C1(new_n464), .C2(new_n463), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n499), .B2(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT71), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT71), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(new_n512), .A3(G62), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n506), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT72), .A3(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n503), .A2(KEYINPUT6), .A3(new_n504), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n509), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n521), .A2(G543), .A3(new_n519), .A4(new_n517), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n514), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n509), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n524), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(G51), .B2(new_n535), .ZN(G168));
  INV_X1    g111(.A(new_n522), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n506), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n537), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n535), .A2(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n506), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  AND3_X1   g129(.A1(new_n521), .A2(new_n519), .A3(new_n517), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n555), .A2(new_n556), .A3(G53), .A4(G543), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n524), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n507), .A2(new_n508), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n537), .A2(G91), .B1(G651), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  XNOR2_X1  g142(.A(G168), .B(new_n567), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G49), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI221_X1 g147(.A(new_n570), .B1(new_n524), .B2(new_n571), .C1(new_n522), .C2(new_n572), .ZN(G288));
  NAND4_X1  g148(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n520), .A2(G86), .A3(new_n509), .A4(new_n521), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n507), .B2(new_n508), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n505), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(G305));
  NAND2_X1  g156(.A1(new_n537), .A2(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n535), .A2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n506), .C2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n587));
  NAND3_X1  g162(.A1(new_n537), .A2(G92), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n535), .A2(G54), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n516), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n587), .B1(new_n537), .B2(G92), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n586), .B1(new_n593), .B2(G868), .ZN(G321));
  XOR2_X1   g169(.A(G321), .B(KEYINPUT77), .Z(G284));
  NOR2_X1   g170(.A1(G299), .A2(G868), .ZN(new_n596));
  XNOR2_X1  g171(.A(G168), .B(KEYINPUT74), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  AOI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  XNOR2_X1  g174(.A(KEYINPUT78), .B(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(G860), .B2(new_n600), .ZN(G148));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n548), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n593), .A2(new_n600), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n484), .A2(G123), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n462), .A2(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  INV_X1    g184(.A(G135), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n607), .B1(new_n608), .B2(new_n609), .C1(new_n610), .C2(new_n487), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND3_X1  g187(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g190(.A(G2100), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n612), .A2(new_n617), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n633), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(G401));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT17), .Z(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n637), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(KEYINPUT81), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(KEYINPUT81), .B2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n639), .A3(new_n637), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n638), .A2(new_n642), .A3(new_n640), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2096), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1991), .B(G1996), .Z(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n664));
  OR2_X1    g239(.A1(new_n662), .A2(new_n660), .ZN(new_n665));
  OAI221_X1 g240(.A(new_n661), .B1(new_n663), .B2(new_n664), .C1(new_n665), .C2(new_n657), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OR3_X1    g242(.A1(new_n666), .A2(KEYINPUT83), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(KEYINPUT83), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n668), .B2(new_n669), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n654), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n673), .ZN(new_n675));
  INV_X1    g250(.A(new_n654), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n676), .A3(new_n671), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  AND3_X1   g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  MUX2_X1   g256(.A(G24), .B(G290), .S(G16), .Z(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G1986), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n484), .A2(G119), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n462), .A2(G107), .ZN(new_n685));
  OAI21_X1  g260(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n686));
  INV_X1    g261(.A(G131), .ZN(new_n687));
  OAI221_X1 g262(.A(new_n684), .B1(new_n685), .B2(new_n686), .C1(new_n687), .C2(new_n487), .ZN(new_n688));
  MUX2_X1   g263(.A(G25), .B(new_n688), .S(G29), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT35), .B(G1991), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G6), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT75), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n580), .B(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n693), .B1(new_n695), .B2(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n692), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n692), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n696), .A2(new_n697), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n698), .A2(new_n703), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n683), .B(new_n691), .C1(new_n709), .C2(KEYINPUT34), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT84), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT85), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(KEYINPUT36), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT93), .B(G1956), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n692), .A2(G20), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G299), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n692), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n719), .A2(G2090), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n692), .A2(G4), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n593), .B2(new_n692), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT86), .B(G1348), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n692), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n549), .B2(new_n692), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1341), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n726), .A2(new_n720), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n727), .B(new_n737), .C1(G2090), .C2(new_n719), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n692), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n692), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT89), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n716), .B1(new_n743), .B2(G34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT88), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT88), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n743), .B2(G34), .ZN(new_n747));
  AOI22_X1  g322(.A1(G160), .A2(G29), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2084), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n716), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n488), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n484), .A2(G128), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(new_n716), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT30), .B(G28), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n761), .A2(new_n716), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n611), .B2(new_n716), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n766));
  NAND3_X1  g341(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G139), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n768), .B1(new_n769), .B2(new_n487), .C1(new_n462), .C2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G29), .B2(G33), .ZN(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n765), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n716), .A2(G32), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n484), .A2(G129), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n782));
  INV_X1    g357(.A(G141), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n487), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n777), .B1(new_n785), .B2(new_n716), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AND4_X1   g363(.A1(new_n749), .A2(new_n760), .A3(new_n776), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G164), .A2(new_n716), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G27), .B2(new_n716), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n793), .B(new_n794), .C1(new_n774), .C2(new_n775), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G1966), .B2(new_n740), .ZN(new_n796));
  NOR2_X1   g371(.A1(G5), .A2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT90), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G301), .B2(new_n692), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1961), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n789), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n738), .A2(new_n742), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n714), .B2(KEYINPUT36), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n715), .A2(new_n803), .ZN(G311));
  INV_X1    g379(.A(G311), .ZN(G150));
  NAND2_X1  g380(.A1(new_n593), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT38), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n522), .A2(new_n808), .B1(new_n524), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n812), .A2(new_n813), .B1(new_n506), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(new_n548), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n548), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n807), .B(new_n818), .Z(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n820), .A2(new_n821), .A3(G860), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n815), .A2(G860), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n479), .B(new_n611), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G162), .Z(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n484), .A2(G126), .B1(new_n492), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n462), .A2(G138), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n467), .B2(new_n468), .ZN(new_n832));
  INV_X1    g407(.A(new_n500), .ZN(new_n833));
  NOR2_X1   g408(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n501), .B(KEYINPUT95), .C1(new_n832), .C2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(KEYINPUT95), .B1(new_n499), .B2(new_n501), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n830), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n757), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n501), .B1(new_n832), .B2(new_n835), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n494), .B1(new_n843), .B2(new_n836), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n756), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n785), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n840), .A2(new_n845), .A3(new_n785), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT96), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n771), .B1(new_n850), .B2(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n484), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n462), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G142), .B2(new_n488), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n614), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n688), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  INV_X1    g436(.A(new_n849), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n785), .B1(new_n840), .B2(new_n845), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT97), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n848), .A2(new_n865), .A3(new_n849), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n861), .B1(new_n867), .B2(new_n771), .ZN(new_n868));
  AOI211_X1 g443(.A(KEYINPUT98), .B(new_n772), .C1(new_n864), .C2(new_n866), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n853), .B(new_n860), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT99), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n862), .A2(KEYINPUT97), .A3(new_n863), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n865), .B1(new_n848), .B2(new_n849), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n771), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT98), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n861), .A3(new_n771), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n875), .A2(new_n876), .B1(new_n851), .B2(new_n852), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT100), .B1(new_n877), .B2(new_n860), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n853), .B1(new_n868), .B2(new_n869), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n880));
  INV_X1    g455(.A(new_n860), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n827), .B1(new_n871), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n870), .B(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n827), .B1(new_n879), .B2(new_n881), .ZN(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n884), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(G395));
  OR2_X1    g467(.A1(new_n591), .A2(new_n592), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n725), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n593), .A2(G299), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT102), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n818), .B(new_n604), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n894), .A2(new_n895), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(G305), .B(G290), .ZN(new_n910));
  XNOR2_X1  g485(.A(G166), .B(G288), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n904), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n909), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n914), .B1(new_n909), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n815), .A2(new_n602), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NOR2_X1   g498(.A1(G286), .A2(G301), .ZN(new_n924));
  NOR2_X1   g499(.A1(G171), .A2(G168), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n817), .B(new_n816), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n597), .B2(G171), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n818), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n906), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n902), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n914), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n912), .B2(new_n913), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n905), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n930), .B1(new_n896), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n940), .B2(new_n929), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(new_n929), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n900), .B1(new_n939), .B2(new_n896), .ZN(new_n945));
  INV_X1    g520(.A(new_n901), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n947), .B2(new_n930), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n937), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n933), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n923), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n933), .B2(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n914), .B(new_n944), .C1(new_n947), .C2(new_n930), .ZN(new_n955));
  AND4_X1   g530(.A1(new_n954), .A2(new_n941), .A3(new_n955), .A4(new_n950), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n953), .A2(new_n956), .A3(KEYINPUT44), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n952), .A2(new_n957), .ZN(G397));
  NAND4_X1  g533(.A1(new_n472), .A2(G40), .A3(new_n478), .A4(new_n473), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n843), .A2(new_n836), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n960), .B2(new_n830), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n830), .B2(new_n841), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT105), .B1(new_n964), .B2(new_n962), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n731), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n959), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n839), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G2067), .ZN(new_n973));
  NOR4_X1   g548(.A1(new_n969), .A2(KEYINPUT60), .A3(new_n893), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n593), .B1(new_n969), .B2(new_n973), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n839), .A2(new_n962), .A3(new_n971), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n970), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n730), .ZN(new_n978));
  INV_X1    g553(.A(new_n973), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n893), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n974), .B1(new_n981), .B2(KEYINPUT60), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n839), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n830), .A2(new_n841), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n971), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n959), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT58), .B(G1341), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n972), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n549), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT116), .B1(new_n993), .B2(KEYINPUT59), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n548), .B1(new_n989), .B2(new_n991), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT59), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND4_X1   g573(.A1(KEYINPUT117), .A2(new_n992), .A3(new_n997), .A4(new_n549), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT117), .B1(new_n995), .B2(new_n997), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n994), .A2(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n982), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n983), .A2(new_n987), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT56), .B(G2072), .Z(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT114), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT50), .B1(new_n844), .B2(G1384), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n959), .B1(new_n962), .B2(new_n964), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1956), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT109), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1012), .B(G1956), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n560), .A2(KEYINPUT110), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n557), .A2(new_n1018), .A3(new_n559), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n565), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1024), .A3(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n560), .A2(new_n565), .A3(KEYINPUT57), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT112), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1016), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n564), .A2(G651), .ZN(new_n1030));
  INV_X1    g605(.A(G91), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n522), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n560), .B2(KEYINPUT110), .ZN(new_n1033));
  AOI211_X1 g608(.A(KEYINPUT111), .B(KEYINPUT57), .C1(new_n1033), .C2(new_n1019), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1024), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1028), .B(new_n1016), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1015), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT61), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1028), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1014), .B1(new_n1042), .B2(new_n1036), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT61), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1002), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1036), .A3(new_n1014), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n975), .B(KEYINPUT115), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT118), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1046), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1047), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n1038), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1042), .A2(new_n1036), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT61), .B1(new_n1054), .B2(new_n1015), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1039), .B(new_n1014), .C1(new_n1042), .C2(new_n1036), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1052), .B(new_n1053), .C1(new_n1057), .C2(new_n1002), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n983), .A2(new_n987), .A3(new_n792), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT120), .B(G1961), .Z(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1065), .B1(new_n977), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT45), .B1(new_n839), .B2(new_n971), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n478), .B1(new_n985), .B2(new_n986), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n474), .A2(G40), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n983), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n986), .B1(new_n844), .B2(G1384), .ZN(new_n1076));
  OR3_X1    g651(.A1(new_n476), .A2(KEYINPUT122), .A3(new_n477), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT122), .B1(new_n476), .B2(new_n477), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(G2105), .A3(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1076), .A2(G40), .A3(new_n474), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1070), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1076), .A2(KEYINPUT123), .A3(new_n1083), .A4(new_n1079), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(KEYINPUT124), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1087), .B(new_n1075), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1067), .B(G301), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1059), .B1(new_n1074), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n977), .A2(new_n1066), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1065), .ZN(new_n1092));
  OAI211_X1 g667(.A(G301), .B(new_n1091), .C1(new_n1092), .C2(new_n1063), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1072), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1067), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n972), .A2(G8), .ZN(new_n1098));
  INV_X1    g673(.A(G1976), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G288), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT52), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1981), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n574), .A2(new_n575), .A3(new_n1102), .A4(new_n579), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT106), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n580), .A2(new_n1106), .A3(G1981), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n580), .B2(G1981), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n961), .B2(new_n970), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n580), .A2(G1981), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT49), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n580), .A2(new_n1106), .A3(G1981), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1104), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1100), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT52), .B1(G288), .B2(new_n1099), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1101), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G166), .A2(new_n1110), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT55), .ZN(new_n1122));
  INV_X1    g697(.A(G2090), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n963), .A2(new_n1123), .A3(new_n968), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1003), .A2(new_n706), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1110), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1120), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT107), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1008), .A2(new_n1123), .A3(new_n1009), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1971), .B1(new_n983), .B2(new_n987), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1008), .A2(new_n1123), .A3(new_n1009), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1125), .A2(KEYINPUT107), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1133), .A3(G8), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1122), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1071), .A2(G1966), .B1(new_n977), .B2(G2084), .ZN(new_n1137));
  INV_X1    g712(.A(G168), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(G8), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(G8), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(KEYINPUT51), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n1142));
  OAI221_X1 g717(.A(G168), .B1(new_n977), .B2(G2084), .C1(new_n1071), .C2(G1966), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(G8), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1127), .B(new_n1136), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1090), .A2(new_n1097), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1049), .A2(new_n1058), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1074), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT62), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1110), .B1(new_n1150), .B2(new_n1128), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1122), .B1(new_n1151), .B2(new_n1133), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(new_n1122), .A3(G8), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1101), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1140), .A2(KEYINPUT51), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1143), .A2(new_n1142), .A3(G8), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1139), .ZN(new_n1161));
  AND4_X1   g736(.A1(new_n1148), .A2(new_n1149), .A3(new_n1157), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT108), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1154), .A2(new_n1120), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1116), .A2(new_n1099), .A3(new_n700), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1103), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1111), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1137), .A2(G8), .A3(new_n597), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1127), .A2(new_n1136), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1126), .A2(new_n1122), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1137), .A2(KEYINPUT63), .A3(G8), .A4(new_n597), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1156), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1163), .B(new_n1167), .C1(new_n1171), .C2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1169), .A2(new_n1170), .B1(new_n1127), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1167), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT108), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1162), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1147), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1076), .A2(new_n959), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n756), .B(new_n759), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n785), .B(G1996), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n688), .B(new_n690), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G290), .B(G1986), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1182), .ZN(new_n1191));
  INV_X1    g766(.A(new_n690), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n688), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1185), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n757), .A2(new_n759), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1191), .A2(G1986), .A3(G290), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT48), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1197), .A2(new_n1198), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1191), .B2(G1996), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1182), .A2(KEYINPUT46), .A3(new_n988), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1183), .A2(new_n785), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1203), .B(new_n1204), .C1(new_n1191), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT47), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1201), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT125), .Z(new_n1211));
  NAND2_X1  g786(.A1(new_n1190), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g787(.A(G319), .ZN(new_n1214));
  NOR3_X1   g788(.A1(G401), .A2(G227), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n1215), .B1(new_n679), .B2(new_n680), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(KEYINPUT126), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1218));
  OAI211_X1 g792(.A(new_n1218), .B(new_n1215), .C1(new_n679), .C2(new_n680), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1220), .B1(new_n953), .B2(new_n956), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1221), .B1(new_n884), .B2(new_n888), .ZN(G308));
  NAND2_X1  g796(.A1(new_n884), .A2(new_n888), .ZN(new_n1223));
  OAI211_X1 g797(.A(new_n1223), .B(new_n1220), .C1(new_n953), .C2(new_n956), .ZN(G225));
endmodule


