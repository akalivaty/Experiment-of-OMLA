//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G77), .ZN(new_n208));
  AND2_X1   g0008(.A1(new_n208), .A2(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G58), .A2(G232), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n207), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n207), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G87), .B(G97), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n220), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n221), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n245), .A2(G20), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n243), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(G50), .B1(new_n221), .B2(G1), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n259), .A2(new_n260), .B1(G50), .B2(new_n256), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g0062(.A(new_n262), .B(KEYINPUT9), .Z(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1698), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(new_n208), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n267), .B(new_n269), .C1(new_n270), .C2(new_n268), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n220), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(G274), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n275), .B2(new_n276), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT66), .A3(new_n282), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n282), .B1(new_n275), .B2(new_n276), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G226), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n279), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n263), .B1(KEYINPUT69), .B2(new_n294), .C1(new_n295), .C2(new_n293), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(KEYINPUT69), .B2(new_n294), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT16), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT7), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n268), .B2(G20), .ZN(new_n302));
  AND2_X1   g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  NOR2_X1   g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n202), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G58), .A2(G68), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n221), .B1(new_n203), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G159), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n246), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n300), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(KEYINPUT74), .B(new_n300), .C1(new_n307), .C2(new_n312), .ZN(new_n316));
  INV_X1    g0116(.A(new_n306), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n305), .B2(new_n221), .ZN(new_n318));
  OAI21_X1  g0118(.A(G68), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT73), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n309), .A2(new_n311), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n309), .B2(new_n311), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n319), .A2(KEYINPUT16), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n315), .A2(new_n243), .A3(new_n316), .A4(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n249), .B1(new_n255), .B2(G20), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n258), .B1(new_n257), .B2(new_n249), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  INV_X1    g0128(.A(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G226), .B2(new_n329), .ZN(new_n331));
  INV_X1    g0131(.A(G87), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n331), .A2(new_n305), .B1(new_n245), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n278), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n291), .A2(G232), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n290), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G169), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n336), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT18), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n336), .A2(new_n295), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(G200), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(new_n326), .A3(new_n324), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n327), .A2(new_n348), .A3(new_n339), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n344), .A2(KEYINPUT17), .A3(new_n326), .A4(new_n324), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n341), .A2(new_n347), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n262), .B1(new_n293), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(G179), .B2(new_n293), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G107), .ZN(new_n357));
  INV_X1    g0157(.A(new_n266), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n356), .B1(new_n357), .B2(new_n268), .C1(new_n358), .C2(new_n227), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n278), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n286), .A2(new_n289), .B1(G244), .B2(new_n291), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  OAI21_X1  g0163(.A(G77), .B1(new_n221), .B2(G1), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n259), .A2(new_n364), .B1(new_n208), .B2(new_n256), .ZN(new_n365));
  INV_X1    g0165(.A(new_n246), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n250), .A2(new_n366), .B1(new_n208), .B2(G20), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT68), .ZN(new_n369));
  INV_X1    g0169(.A(new_n251), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n365), .B1(new_n371), .B2(new_n243), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n363), .B(new_n372), .C1(new_n295), .C2(new_n362), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(new_n362), .B2(new_n353), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n360), .A2(new_n338), .A3(new_n361), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n299), .A2(new_n352), .A3(new_n355), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT70), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n284), .A2(new_n285), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT66), .B1(new_n288), .B2(new_n282), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n227), .A2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G226), .B2(G1698), .ZN(new_n385));
  INV_X1    g0185(.A(G97), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n385), .A2(new_n305), .B1(new_n245), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n278), .B1(new_n291), .B2(G238), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT71), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n379), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n383), .A2(new_n388), .A3(KEYINPUT71), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n383), .A2(new_n388), .A3(new_n379), .A4(new_n389), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(G179), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n395), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT14), .B1(new_n398), .B2(G169), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n400), .B(new_n353), .C1(new_n397), .C2(new_n395), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n251), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n403));
  INV_X1    g0203(.A(G50), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n246), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT11), .B1(new_n405), .B2(new_n243), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT72), .B1(new_n256), .B2(G68), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT12), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(KEYINPUT11), .A3(new_n243), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n258), .B(G68), .C1(G1), .C2(new_n221), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n394), .A2(G190), .A3(new_n395), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n398), .B2(G200), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n402), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n378), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G283), .ZN(new_n418));
  OAI211_X1 g0218(.A(G250), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n419));
  OAI211_X1 g0219(.A(G244), .B(new_n329), .C1(new_n303), .C2(new_n304), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT4), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT4), .B1(new_n266), .B2(G244), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n278), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT5), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G41), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n280), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(KEYINPUT77), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n280), .A2(KEYINPUT5), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n255), .A2(G45), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n288), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT77), .B1(new_n427), .B2(new_n428), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n281), .A2(G1), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n426), .A2(G41), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n427), .A2(new_n428), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G257), .A3(new_n283), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n424), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n433), .B2(new_n435), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n424), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(G190), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT79), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n444), .A2(KEYINPUT79), .A3(G190), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n442), .A2(G200), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n257), .A2(new_n386), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n255), .A2(G33), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n244), .A2(new_n256), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n453), .B1(new_n456), .B2(new_n386), .ZN(new_n457));
  OAI21_X1  g0257(.A(G107), .B1(new_n317), .B2(new_n318), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n366), .A2(G77), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT6), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(KEYINPUT6), .B2(new_n386), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT75), .B(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n458), .B(new_n459), .C1(new_n464), .C2(new_n221), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n457), .B1(new_n465), .B2(new_n243), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n221), .B(G87), .C1(new_n303), .C2(new_n304), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT22), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n268), .A2(new_n470), .A3(new_n221), .A4(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n357), .A2(G20), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT23), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n473), .B2(KEYINPUT23), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n473), .B2(KEYINPUT23), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n472), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n472), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n243), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT84), .B(new_n243), .C1(new_n482), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n440), .A2(G264), .A3(new_n283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT85), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT85), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n440), .A2(new_n491), .A3(G264), .A4(new_n283), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G294), .ZN(new_n495));
  INV_X1    g0295(.A(G250), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n495), .C1(new_n358), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n278), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n498), .A3(new_n437), .ZN(new_n499));
  INV_X1    g0299(.A(G200), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n490), .A2(new_n492), .B1(new_n497), .B2(new_n278), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n295), .A3(new_n437), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT86), .ZN(new_n504));
  OR3_X1    g0304(.A1(new_n499), .A2(KEYINPUT86), .A3(G190), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n357), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT25), .B1(new_n257), .B2(new_n357), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n456), .A2(new_n357), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n488), .A2(new_n504), .A3(new_n505), .A4(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n442), .A2(G179), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n466), .A2(new_n512), .ZN(new_n513));
  AND4_X1   g0313(.A1(KEYINPUT78), .A2(new_n424), .A3(new_n437), .A4(new_n441), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT78), .B1(new_n446), .B2(new_n424), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n353), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n467), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n488), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n499), .A2(new_n353), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(G179), .B2(new_n499), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G244), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n524));
  OAI211_X1 g0324(.A(G238), .B(new_n329), .C1(new_n303), .C2(new_n304), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n278), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n496), .B1(new_n281), .B2(G1), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n255), .A2(new_n287), .A3(G45), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n283), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT80), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n534), .B(new_n531), .C1(new_n527), .C2(new_n278), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n338), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n370), .B2(new_n386), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n268), .A2(new_n221), .A3(G68), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g0341(.A(KEYINPUT81), .B(G87), .Z(new_n542));
  NAND3_X1  g0342(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n460), .B1(new_n221), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n243), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n369), .A2(new_n257), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n369), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n455), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n353), .B1(new_n533), .B2(new_n535), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n537), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n536), .A2(G190), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n545), .B(new_n546), .C1(new_n332), .C2(new_n456), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n533), .B2(new_n535), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n427), .A2(new_n428), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n438), .A2(new_n439), .ZN(new_n562));
  OAI211_X1 g0362(.A(G270), .B(new_n283), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT82), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n440), .A2(KEYINPUT82), .A3(G270), .A4(new_n283), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G264), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(new_n329), .C1(new_n303), .C2(new_n304), .ZN(new_n569));
  INV_X1    g0369(.A(G303), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n268), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n278), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n567), .A2(new_n437), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n418), .B(new_n221), .C1(G33), .C2(new_n386), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n243), .C1(new_n221), .C2(G116), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n256), .A2(G116), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n455), .B2(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(G169), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n573), .A2(G200), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n565), .A2(new_n566), .B1(new_n434), .B2(new_n436), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G190), .A3(new_n572), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n338), .B1(new_n571), .B2(new_n278), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n580), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n573), .A2(new_n580), .A3(KEYINPUT21), .A4(G169), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n583), .A2(new_n588), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n523), .A2(new_n560), .A3(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n417), .A2(new_n518), .A3(new_n593), .ZN(G372));
  INV_X1    g0394(.A(new_n349), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n348), .B1(new_n327), .B2(new_n339), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n347), .A2(new_n350), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n402), .A2(new_n412), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n413), .A2(new_n414), .ZN(new_n602));
  INV_X1    g0402(.A(new_n376), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n299), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(new_n355), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n536), .A2(new_n338), .B1(new_n548), .B2(new_n550), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n528), .A2(new_n532), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n353), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n555), .B1(new_n536), .B2(G190), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n500), .B1(new_n528), .B2(new_n532), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT87), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n608), .A2(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n467), .A2(new_n511), .A3(new_n614), .A4(new_n517), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n509), .B1(new_n486), .B2(new_n487), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n521), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT26), .B1(new_n559), .B2(new_n517), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n537), .A2(new_n551), .A3(new_n610), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n611), .A2(new_n613), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(new_n622), .A3(new_n513), .A4(new_n516), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n621), .B(new_n622), .C1(KEYINPUT26), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n607), .B1(new_n417), .B2(new_n626), .ZN(G369));
  NAND3_X1  g0427(.A1(new_n255), .A2(new_n221), .A3(G13), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT88), .ZN(new_n630));
  INV_X1    g0430(.A(G213), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n628), .B2(KEYINPUT27), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT89), .A3(G343), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n585), .ZN(new_n641));
  MUX2_X1   g0441(.A(new_n592), .B(new_n618), .S(new_n641), .Z(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n523), .A2(new_n639), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n511), .B1(new_n616), .B2(new_n640), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n523), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n639), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(G399));
  INV_X1    g0452(.A(new_n217), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G41), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n224), .ZN(new_n655));
  INV_X1    g0455(.A(G116), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n542), .A2(new_n656), .A3(new_n460), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G1), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  AOI21_X1  g0460(.A(G179), .B1(new_n528), .B2(new_n532), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n499), .A2(new_n573), .A3(new_n442), .A4(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n514), .A2(new_n515), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n493), .A2(new_n498), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n665), .A2(new_n533), .A3(new_n535), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n567), .A2(new_n437), .A3(new_n589), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT90), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n586), .A2(new_n669), .A3(new_n589), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n664), .A2(new_n666), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT92), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n444), .A2(new_n447), .A3(new_n536), .A4(new_n502), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n670), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT92), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(KEYINPUT30), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n663), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT30), .B1(new_n671), .B2(KEYINPUT91), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n669), .A2(new_n567), .A3(new_n437), .A4(new_n589), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n669), .B1(new_n586), .B2(new_n589), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT91), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(new_n664), .A4(new_n666), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT93), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT91), .B1(new_n674), .B2(new_n675), .ZN(new_n687));
  AND4_X1   g0487(.A1(KEYINPUT93), .A2(new_n685), .A3(new_n687), .A4(new_n672), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n679), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT31), .B1(new_n689), .B2(new_n639), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n467), .A2(new_n511), .A3(new_n517), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n617), .A2(new_n559), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n592), .A3(new_n692), .A4(new_n640), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n685), .A2(new_n687), .A3(new_n672), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n677), .B1(new_n676), .B2(KEYINPUT30), .ZN(new_n695));
  NOR4_X1   g0495(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT92), .A4(new_n672), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n694), .B(new_n662), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n640), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n693), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n690), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT95), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n617), .B2(new_n618), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n649), .B(KEYINPUT95), .C1(new_n616), .C2(new_n521), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n622), .B1(new_n708), .B2(new_n615), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT26), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n624), .A2(KEYINPUT94), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n559), .B2(new_n517), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n624), .A2(new_n710), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(KEYINPUT29), .B(new_n640), .C1(new_n709), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n626), .A2(new_n639), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(KEYINPUT29), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n704), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n660), .B1(new_n720), .B2(G1), .ZN(G364));
  INV_X1    g0521(.A(G13), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n255), .B1(new_n723), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n654), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n644), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G330), .B2(new_n642), .ZN(new_n728));
  INV_X1    g0528(.A(new_n726), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n220), .B1(G20), .B2(new_n353), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n221), .ZN(new_n733));
  INV_X1    g0533(.A(G294), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n221), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n295), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(G283), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n733), .A2(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n295), .A3(new_n500), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n268), .B1(new_n740), .B2(G329), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n570), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n295), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n738), .B(new_n743), .C1(G326), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(G190), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT33), .B(G317), .ZN(new_n749));
  NAND2_X1  g0549(.A1(G20), .A2(G179), .ZN(new_n750));
  AOI21_X1  g0550(.A(G200), .B1(new_n750), .B2(KEYINPUT96), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(KEYINPUT96), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n295), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n748), .A2(new_n749), .B1(new_n753), .B2(G322), .ZN(new_n754));
  INV_X1    g0554(.A(G311), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n747), .B(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n733), .A2(new_n386), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n542), .A2(new_n742), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n736), .A2(new_n357), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n305), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G50), .A2(new_n746), .B1(new_n748), .B2(G68), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G58), .A2(new_n753), .B1(new_n756), .B2(new_n208), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n739), .A2(new_n310), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n731), .B1(new_n758), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n730), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n217), .A2(G355), .A3(new_n268), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n653), .A2(new_n268), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G45), .B2(new_n223), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n240), .A2(G45), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n773), .B1(G116), .B2(new_n217), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n729), .B(new_n768), .C1(new_n772), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n771), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n642), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n728), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(G396));
  OR2_X1    g0582(.A1(new_n640), .A2(new_n372), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n603), .B1(new_n783), .B2(new_n373), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n376), .A2(new_n639), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n718), .B(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n726), .B1(new_n787), .B2(new_n704), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n704), .B2(new_n787), .ZN(new_n789));
  INV_X1    g0589(.A(G77), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n730), .A2(new_n769), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n729), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n268), .B(new_n759), .C1(G311), .C2(new_n740), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n736), .A2(new_n332), .ZN(new_n794));
  INV_X1    g0594(.A(new_n742), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G107), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n753), .ZN(new_n798));
  INV_X1    g0598(.A(new_n746), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n734), .B2(new_n798), .C1(new_n570), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n748), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n801), .A2(new_n737), .B1(new_n757), .B2(new_n656), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(KEYINPUT98), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(KEYINPUT98), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G143), .A2(new_n753), .B1(new_n756), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n806), .B2(new_n799), .C1(new_n247), .C2(new_n801), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT34), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n736), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G68), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n268), .C1(new_n812), .C2(new_n739), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n733), .A2(new_n201), .B1(new_n742), .B2(new_n404), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n807), .C2(new_n808), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n803), .A2(new_n804), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n792), .B1(new_n816), .B2(new_n731), .C1(new_n770), .C2(new_n786), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n789), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G384));
  NOR2_X1   g0619(.A1(new_n723), .A2(new_n255), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n321), .A2(new_n322), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n300), .B1(new_n821), .B2(new_n307), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n243), .A3(new_n323), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n823), .A2(new_n824), .A3(new_n326), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n823), .B2(new_n326), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n339), .A2(new_n634), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n345), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT37), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n327), .A2(new_n634), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n340), .A2(new_n831), .A3(new_n345), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n825), .A2(new_n826), .A3(new_n633), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n351), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT38), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT38), .B1(new_n834), .B2(new_n836), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT39), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n340), .A2(new_n831), .A3(new_n345), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n833), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n831), .B1(new_n599), .B2(new_n597), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT39), .B1(new_n848), .B2(new_n837), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n402), .A2(new_n412), .A3(new_n640), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n838), .A2(new_n839), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n640), .B(new_n786), .C1(new_n620), .C2(new_n625), .ZN(new_n856));
  INV_X1    g0656(.A(new_n785), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n398), .A2(G169), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n400), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n398), .A2(KEYINPUT14), .A3(G169), .ZN(new_n860));
  INV_X1    g0660(.A(new_n395), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n392), .B2(new_n393), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n859), .A2(new_n860), .B1(G179), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n602), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n639), .A2(new_n412), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n865), .B1(new_n863), .B2(new_n602), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n870), .A2(KEYINPUT100), .B1(new_n415), .B2(new_n865), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n856), .A2(new_n857), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n855), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n598), .A2(new_n633), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n853), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n607), .B1(new_n417), .B2(new_n719), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n875), .B(new_n876), .Z(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n601), .A2(new_n602), .A3(new_n865), .ZN(new_n879));
  INV_X1    g0679(.A(new_n602), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT100), .B(new_n866), .C1(new_n880), .C2(new_n402), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT100), .B1(new_n864), .B2(new_n866), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n786), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n662), .B1(new_n695), .B2(new_n696), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT93), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n694), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n680), .A2(KEYINPUT93), .A3(new_n685), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n699), .B1(new_n889), .B2(new_n640), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n593), .A2(new_n518), .A3(new_n639), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n689), .B2(new_n700), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n884), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n855), .B1(new_n893), .B2(KEYINPUT102), .ZN(new_n894));
  INV_X1    g0694(.A(new_n786), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n871), .B2(new_n869), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n693), .B1(new_n889), .B2(new_n701), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n690), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n878), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n351), .A2(new_n327), .A3(new_n634), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n902), .B2(new_n845), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT40), .B1(new_n838), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n893), .B2(KEYINPUT103), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n897), .A2(new_n690), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n909), .B1(new_n417), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n378), .A2(new_n416), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n890), .A2(new_n892), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n901), .A2(new_n912), .A3(new_n913), .A4(new_n908), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(G330), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n820), .B1(new_n877), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n877), .B2(new_n915), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT35), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n464), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n464), .A2(new_n918), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(G116), .A3(new_n222), .A4(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n224), .A2(new_n208), .A3(new_n308), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(G50), .B2(new_n202), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n722), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT99), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n917), .A2(new_n927), .ZN(G367));
  NOR2_X1   g0728(.A1(new_n517), .A2(new_n640), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT104), .Z(new_n930));
  OAI211_X1 g0730(.A(new_n467), .B(new_n517), .C1(new_n466), .C2(new_n640), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n647), .A3(new_n650), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n934), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n932), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n517), .B1(new_n937), .B2(new_n523), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n938), .A2(new_n640), .B1(KEYINPUT42), .B2(new_n933), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n639), .A2(new_n555), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n614), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n622), .B2(new_n941), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT43), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(KEYINPUT106), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n936), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT106), .B1(new_n940), .B2(new_n944), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n948), .A2(new_n949), .B1(new_n648), .B2(new_n937), .ZN(new_n950));
  INV_X1    g0750(.A(new_n949), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n648), .A2(new_n937), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n947), .A4(new_n945), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n654), .B(KEYINPUT41), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n651), .A2(new_n932), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT45), .Z(new_n956));
  NOR2_X1   g0756(.A1(new_n651), .A2(new_n932), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n648), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n647), .B(new_n650), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT107), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(new_n643), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n643), .B(KEYINPUT107), .Z(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n956), .A2(new_n648), .A3(new_n958), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n961), .A2(new_n720), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n954), .B1(new_n968), .B2(new_n720), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n950), .B(new_n953), .C1(new_n969), .C2(new_n725), .ZN(new_n970));
  INV_X1    g0770(.A(new_n774), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n772), .B1(new_n217), .B2(new_n369), .C1(new_n971), .C2(new_n233), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n726), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n801), .A2(new_n310), .ZN(new_n974));
  XNOR2_X1  g0774(.A(KEYINPUT109), .B(G137), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n268), .B1(new_n739), .B2(new_n975), .C1(new_n733), .C2(new_n202), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n270), .A2(new_n736), .B1(new_n742), .B2(new_n201), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n746), .A2(G143), .B1(new_n753), .B2(G150), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n404), .C2(new_n757), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n734), .A2(new_n801), .B1(new_n799), .B2(new_n755), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G303), .B2(new_n753), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n268), .B1(new_n740), .B2(G317), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n386), .B2(new_n736), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n795), .A2(G116), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n982), .B(new_n987), .C1(new_n985), .C2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(new_n733), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n756), .A2(G283), .B1(G107), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT108), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n980), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n973), .B1(new_n779), .B2(new_n943), .C1(new_n993), .C2(new_n731), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n970), .A2(new_n994), .ZN(G387));
  NOR2_X1   g0795(.A1(new_n966), .A2(new_n720), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT112), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n966), .A2(new_n720), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n654), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n966), .A2(new_n725), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n230), .A2(new_n281), .A3(new_n268), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT50), .B1(new_n249), .B2(G50), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n281), .C1(new_n202), .C2(new_n790), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n249), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n305), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n657), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n653), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n772), .B1(new_n217), .B2(new_n357), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n726), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n268), .B1(new_n739), .B2(new_n247), .C1(new_n386), .C2(new_n736), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n208), .B2(new_n795), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n369), .A2(new_n733), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n746), .A2(G159), .B1(new_n756), .B2(G68), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n748), .A2(new_n250), .B1(new_n753), .B2(G50), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n733), .A2(new_n737), .B1(new_n742), .B2(new_n734), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G311), .A2(new_n748), .B1(new_n746), .B2(G322), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G303), .A2(new_n756), .B1(new_n753), .B2(G317), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  AOI21_X1  g0827(.A(new_n268), .B1(new_n740), .B2(G326), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n656), .B2(new_n736), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT110), .Z(new_n1030));
  OAI21_X1  g0830(.A(new_n1019), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1012), .B1(new_n1031), .B2(new_n730), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n647), .B2(new_n779), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1003), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1002), .A2(new_n1035), .ZN(G393));
  INV_X1    g0836(.A(KEYINPUT113), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n961), .A2(new_n1037), .A3(new_n967), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n967), .A2(new_n1037), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n724), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n937), .A2(new_n771), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n774), .A2(new_n237), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n772), .B1(new_n217), .B2(new_n386), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n726), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n746), .A2(G317), .B1(new_n753), .B2(G311), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n268), .B(new_n761), .C1(G322), .C2(new_n740), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n989), .A2(G116), .B1(new_n795), .B2(G283), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n734), .B2(new_n757), .C1(new_n570), .C2(new_n801), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n305), .B(new_n794), .C1(G143), .C2(new_n740), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n989), .A2(G77), .B1(new_n795), .B2(G68), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n404), .B2(new_n801), .C1(new_n249), .C2(new_n757), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n746), .A2(G150), .B1(new_n753), .B2(G159), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1046), .A2(new_n1050), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1044), .B1(new_n1057), .B2(new_n730), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1040), .B1(new_n1041), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1038), .A2(new_n998), .A3(new_n1039), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n654), .A3(new_n968), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(G390));
  NAND3_X1  g0862(.A1(new_n913), .A2(G330), .A3(new_n786), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n882), .A2(new_n883), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n784), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n640), .B(new_n1066), .C1(new_n709), .C2(new_n716), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1064), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n703), .A2(G330), .A3(new_n786), .A4(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n857), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  OAI211_X1 g0871(.A(G330), .B(new_n786), .C1(new_n690), .C2(new_n702), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1064), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n896), .B(G330), .C1(new_n897), .C2(new_n690), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n856), .A2(new_n857), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1076), .ZN(new_n1078));
  AOI211_X1 g0878(.A(KEYINPUT114), .B(new_n1078), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1070), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(G330), .ZN(new_n1081));
  NOR4_X1   g0881(.A1(new_n910), .A2(new_n378), .A3(new_n1081), .A4(new_n416), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n876), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1074), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1076), .A2(new_n1068), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n840), .B1(new_n838), .B2(new_n903), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n834), .A2(new_n836), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n842), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1086), .A2(new_n851), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n851), .B1(new_n838), .B2(new_n903), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1067), .A2(new_n857), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n1068), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1085), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n841), .A2(new_n849), .B1(new_n872), .B2(new_n852), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1064), .B1(new_n1067), .B2(new_n857), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1069), .C1(new_n1097), .C2(new_n1092), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1084), .A2(KEYINPUT115), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT115), .B1(new_n1084), .B2(new_n1100), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1084), .ZN(new_n1104));
  AOI211_X1 g0904(.A(G41), .B(new_n653), .C1(new_n1104), .C2(new_n1099), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1099), .A2(new_n725), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n791), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n726), .B1(new_n250), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n733), .A2(new_n310), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n305), .B(new_n1110), .C1(G125), .C2(new_n740), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1111), .B1(new_n404), .B2(new_n736), .C1(new_n1112), .C2(new_n799), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G132), .A2(new_n753), .B1(new_n756), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n742), .A2(new_n247), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(new_n801), .C2(new_n975), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n746), .A2(G283), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n989), .A2(G77), .B1(new_n795), .B2(G87), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n268), .B1(new_n740), .B2(G294), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n811), .A4(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n748), .A2(G107), .B1(new_n753), .B2(G116), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n386), .B2(new_n757), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1113), .A2(new_n1119), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1109), .B1(new_n1126), .B2(new_n730), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n850), .B2(new_n770), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1106), .A2(new_n1107), .A3(new_n1128), .ZN(G378));
  AOI21_X1  g0929(.A(new_n854), .B1(new_n898), .B2(new_n899), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n893), .A2(KEYINPUT102), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT40), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n896), .B(KEYINPUT103), .C1(new_n897), .C2(new_n690), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n878), .B1(new_n848), .B2(new_n837), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT103), .B1(new_n913), .B2(new_n896), .ZN(new_n1136));
  OAI21_X1  g0936(.A(G330), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT117), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1081), .B1(new_n905), .B2(new_n907), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n901), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n262), .A2(new_n633), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT116), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n299), .A2(new_n355), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n299), .B2(new_n355), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1148));
  XOR2_X1   g0948(.A(new_n1147), .B(new_n1148), .Z(new_n1149));
  NAND3_X1  g0949(.A1(new_n1138), .A2(new_n1141), .A3(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1147), .B(new_n1148), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n1140), .A3(new_n901), .A4(new_n1139), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n875), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n876), .A2(new_n1082), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1150), .A2(new_n875), .A3(new_n1152), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1155), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT118), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1155), .A2(new_n1159), .A3(KEYINPUT118), .A4(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1150), .A2(new_n875), .A3(new_n1152), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n875), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1157), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT119), .B1(new_n1168), .B2(KEYINPUT57), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1157), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1155), .A2(new_n1170), .A3(new_n1160), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT119), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n1158), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1165), .A2(new_n654), .A3(new_n1169), .A4(new_n1173), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1166), .A2(new_n1167), .A3(new_n724), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1151), .A2(new_n769), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n726), .B1(G50), .B2(new_n1108), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1112), .A2(new_n798), .B1(new_n757), .B2(new_n806), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n989), .A2(G150), .B1(new_n795), .B2(new_n1115), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n801), .B2(new_n812), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G125), .C2(new_n746), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n810), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n740), .C2(G124), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n549), .A2(new_n756), .B1(new_n753), .B2(G107), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n656), .B2(new_n799), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n801), .A2(new_n386), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n268), .A2(G41), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n737), .B2(new_n739), .C1(new_n202), .C2(new_n733), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n270), .A2(new_n742), .B1(new_n736), .B2(new_n201), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1191), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n404), .C1(G33), .C2(G41), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1187), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1177), .B1(new_n1199), .B2(new_n730), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1175), .B1(new_n1176), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1174), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G375));
  OR2_X1    g1003(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n954), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1084), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT120), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1064), .A2(new_n769), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n799), .A2(new_n812), .B1(new_n798), .B2(new_n975), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G150), .B2(new_n756), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n268), .B1(new_n739), .B2(new_n1112), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n733), .A2(new_n404), .B1(new_n742), .B2(new_n310), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G58), .C2(new_n810), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1210), .B(new_n1213), .C1(new_n801), .C2(new_n1114), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n801), .A2(new_n656), .B1(new_n798), .B2(new_n737), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G294), .B2(new_n746), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n268), .B(new_n1015), .C1(G77), .C2(new_n810), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n795), .B1(new_n740), .B2(G303), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT121), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1218), .A2(new_n1219), .B1(new_n756), .B2(G107), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1216), .A2(new_n1217), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n731), .B1(new_n1214), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n729), .B(new_n1223), .C1(new_n202), .C2(new_n791), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1080), .A2(new_n725), .B1(new_n1208), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1207), .A2(new_n1225), .ZN(G381));
  NAND3_X1  g1026(.A1(new_n1002), .A2(new_n781), .A3(new_n1035), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1059), .A2(new_n818), .A3(new_n1061), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(G378), .A2(G387), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1202), .A2(new_n1229), .A3(new_n1225), .A4(new_n1207), .ZN(G407));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n631), .A2(G343), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1202), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(G407), .A2(G213), .A3(new_n1233), .ZN(G409));
  INV_X1    g1034(.A(KEYINPUT123), .ZN(new_n1235));
  AND3_X1   g1035(.A1(G390), .A2(new_n994), .A3(new_n970), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G390), .B1(new_n994), .B2(new_n970), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1227), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n1235), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1174), .A2(G378), .A3(new_n1201), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1201), .B1(new_n954), .B2(new_n1171), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1231), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1232), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1084), .A2(KEYINPUT60), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1249), .A2(new_n1204), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n654), .B1(new_n1249), .B2(new_n1204), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1225), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(G384), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT62), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1232), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT125), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1258), .B(new_n1232), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1253), .A2(KEYINPUT62), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1254), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1232), .A2(G2897), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT122), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1253), .B(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1244), .B1(new_n1262), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1242), .A2(new_n1270), .A3(new_n1243), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1242), .A2(new_n1273), .A3(new_n1243), .A4(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1248), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1265), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1279), .A2(KEYINPUT63), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1269), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(new_n1245), .A2(KEYINPUT127), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1202), .A2(G378), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1284), .A2(new_n1253), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1253), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1244), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1244), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1244), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1283), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1287), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(G402));
endmodule


