

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743;

  BUF_X1 U371 ( .A(n666), .Z(n351) );
  XNOR2_X1 U372 ( .A(n521), .B(KEYINPUT35), .ZN(n738) );
  OR2_X1 U373 ( .A1(n598), .A2(n574), .ZN(n573) );
  NAND2_X1 U374 ( .A1(n371), .A2(n369), .ZN(n521) );
  NOR2_X1 U375 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U376 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U377 ( .A(n501), .B(n500), .ZN(n666) );
  BUF_X1 U378 ( .A(n641), .Z(n352) );
  XNOR2_X1 U379 ( .A(n558), .B(n559), .ZN(n657) );
  NOR2_X1 U380 ( .A1(n640), .A2(n641), .ZN(n484) );
  XNOR2_X1 U381 ( .A(n423), .B(KEYINPUT1), .ZN(n641) );
  NAND2_X1 U382 ( .A1(n366), .A2(n365), .ZN(n423) );
  XNOR2_X1 U383 ( .A(n488), .B(n350), .ZN(n694) );
  XNOR2_X1 U384 ( .A(n727), .B(G146), .ZN(n488) );
  INV_X1 U385 ( .A(n482), .ZN(n350) );
  XNOR2_X1 U386 ( .A(n446), .B(G128), .ZN(n475) );
  XNOR2_X1 U387 ( .A(G116), .B(G113), .ZN(n493) );
  INV_X1 U388 ( .A(G101), .ZN(n490) );
  XNOR2_X2 U389 ( .A(n513), .B(n512), .ZN(n581) );
  XNOR2_X2 U390 ( .A(n562), .B(KEYINPUT41), .ZN(n417) );
  XNOR2_X1 U391 ( .A(n349), .B(n433), .ZN(n403) );
  NAND2_X1 U392 ( .A1(n743), .A2(n742), .ZN(n349) );
  XNOR2_X1 U393 ( .A(G113), .B(G143), .ZN(n435) );
  NOR2_X1 U394 ( .A1(G902), .A2(n705), .ZN(n458) );
  INV_X1 U395 ( .A(G953), .ZN(n734) );
  XNOR2_X1 U396 ( .A(n673), .B(KEYINPUT2), .ZN(n605) );
  XNOR2_X2 U397 ( .A(KEYINPUT40), .B(n573), .ZN(n742) );
  INV_X1 U398 ( .A(KEYINPUT100), .ZN(n401) );
  NOR2_X1 U399 ( .A1(n405), .A2(n403), .ZN(n596) );
  NAND2_X2 U400 ( .A1(n396), .A2(n394), .ZN(n538) );
  NOR2_X1 U401 ( .A1(n588), .A2(n571), .ZN(n572) );
  AND2_X1 U402 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U403 ( .A1(n393), .A2(n395), .ZN(n394) );
  XNOR2_X1 U404 ( .A(n418), .B(n560), .ZN(n662) );
  XNOR2_X1 U405 ( .A(n402), .B(n401), .ZN(n400) );
  XNOR2_X1 U406 ( .A(n495), .B(n353), .ZN(n503) );
  XNOR2_X1 U407 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U408 ( .A1(n492), .A2(n491), .ZN(n494) );
  NOR2_X1 U409 ( .A1(n640), .A2(n423), .ZN(n564) );
  XNOR2_X2 U410 ( .A(n510), .B(n355), .ZN(n558) );
  OR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n511) );
  XOR2_X1 U412 ( .A(G122), .B(G104), .Z(n502) );
  XNOR2_X1 U413 ( .A(n416), .B(G125), .ZN(n507) );
  INV_X1 U414 ( .A(G146), .ZN(n416) );
  XNOR2_X1 U415 ( .A(n499), .B(n361), .ZN(n565) );
  INV_X1 U416 ( .A(G472), .ZN(n361) );
  NAND2_X1 U417 ( .A1(n657), .A2(n656), .ZN(n418) );
  XNOR2_X1 U418 ( .A(n444), .B(n443), .ZN(n533) );
  XNOR2_X1 U419 ( .A(n507), .B(n415), .ZN(n460) );
  INV_X1 U420 ( .A(KEYINPUT10), .ZN(n415) );
  INV_X1 U421 ( .A(n741), .ZN(n390) );
  OR2_X1 U422 ( .A1(n407), .A2(n739), .ZN(n405) );
  XNOR2_X1 U423 ( .A(n738), .B(KEYINPUT67), .ZN(n424) );
  NOR2_X1 U424 ( .A1(n622), .A2(n391), .ZN(n425) );
  NAND2_X1 U425 ( .A1(n390), .A2(n392), .ZN(n391) );
  XNOR2_X1 U426 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n449) );
  XOR2_X1 U427 ( .A(G107), .B(G122), .Z(n448) );
  XNOR2_X1 U428 ( .A(n506), .B(n354), .ZN(n727) );
  XNOR2_X1 U429 ( .A(n384), .B(G110), .ZN(n504) );
  XNOR2_X1 U430 ( .A(G107), .B(KEYINPUT76), .ZN(n384) );
  XNOR2_X1 U431 ( .A(G137), .B(G140), .ZN(n476) );
  XNOR2_X1 U432 ( .A(n475), .B(n474), .ZN(n506) );
  INV_X1 U433 ( .A(KEYINPUT4), .ZN(n474) );
  NOR2_X1 U434 ( .A1(n522), .A2(n533), .ZN(n561) );
  XNOR2_X1 U435 ( .A(n564), .B(n409), .ZN(n570) );
  NAND2_X1 U436 ( .A1(n428), .A2(n427), .ZN(n431) );
  NOR2_X1 U437 ( .A1(n600), .A2(n647), .ZN(n427) );
  INV_X1 U438 ( .A(n527), .ZN(n428) );
  OR2_X1 U439 ( .A1(n694), .A2(n357), .ZN(n365) );
  AND2_X1 U440 ( .A1(n364), .A2(n367), .ZN(n366) );
  XNOR2_X1 U441 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U442 ( .A(KEYINPUT91), .B(KEYINPUT77), .ZN(n411) );
  XNOR2_X1 U443 ( .A(n413), .B(G110), .ZN(n412) );
  INV_X1 U444 ( .A(KEYINPUT24), .ZN(n413) );
  XNOR2_X1 U445 ( .A(n461), .B(n462), .ZN(n414) );
  XNOR2_X1 U446 ( .A(G119), .B(G128), .ZN(n461) );
  XNOR2_X1 U447 ( .A(KEYINPUT71), .B(KEYINPUT23), .ZN(n462) );
  XNOR2_X1 U448 ( .A(n504), .B(n383), .ZN(n481) );
  XNOR2_X1 U449 ( .A(n476), .B(n477), .ZN(n383) );
  XNOR2_X1 U450 ( .A(G101), .B(G104), .ZN(n477) );
  XNOR2_X1 U451 ( .A(n720), .B(n432), .ZN(n687) );
  XNOR2_X1 U452 ( .A(n506), .B(n509), .ZN(n432) );
  XNOR2_X1 U453 ( .A(n422), .B(n419), .ZN(n509) );
  XNOR2_X1 U454 ( .A(n421), .B(n420), .ZN(n419) );
  XNOR2_X1 U455 ( .A(KEYINPUT33), .B(KEYINPUT88), .ZN(n500) );
  INV_X1 U456 ( .A(n538), .ZN(n375) );
  INV_X1 U457 ( .A(n519), .ZN(n374) );
  XNOR2_X1 U458 ( .A(n442), .B(n441), .ZN(n700) );
  NOR2_X1 U459 ( .A1(G952), .A2(n734), .ZN(n712) );
  AND2_X1 U460 ( .A1(n595), .A2(n587), .ZN(n408) );
  INV_X1 U461 ( .A(n561), .ZN(n659) );
  INV_X1 U462 ( .A(KEYINPUT103), .ZN(n409) );
  INV_X1 U463 ( .A(G469), .ZN(n368) );
  NAND2_X1 U464 ( .A1(n368), .A2(G902), .ZN(n367) );
  XNOR2_X1 U465 ( .A(KEYINPUT17), .B(KEYINPUT89), .ZN(n420) );
  XNOR2_X1 U466 ( .A(KEYINPUT78), .B(KEYINPUT18), .ZN(n421) );
  XNOR2_X1 U467 ( .A(n507), .B(n508), .ZN(n422) );
  XNOR2_X1 U468 ( .A(KEYINPUT15), .B(G902), .ZN(n604) );
  NAND2_X1 U469 ( .A1(n644), .A2(n643), .ZN(n640) );
  NOR2_X1 U470 ( .A1(n517), .A2(n399), .ZN(n395) );
  NAND2_X1 U471 ( .A1(n561), .A2(n643), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n362), .B(n488), .ZN(n607) );
  XNOR2_X1 U473 ( .A(n498), .B(n487), .ZN(n362) );
  AND2_X1 U474 ( .A1(n639), .A2(n387), .ZN(n386) );
  INV_X1 U475 ( .A(n637), .ZN(n387) );
  NAND2_X1 U476 ( .A1(n382), .A2(n426), .ZN(n389) );
  XNOR2_X1 U477 ( .A(n385), .B(n505), .ZN(n720) );
  XNOR2_X1 U478 ( .A(n503), .B(n502), .ZN(n385) );
  XNOR2_X1 U479 ( .A(G116), .B(G134), .ZN(n447) );
  INV_X1 U480 ( .A(G143), .ZN(n446) );
  XNOR2_X1 U481 ( .A(G131), .B(G140), .ZN(n436) );
  XOR2_X1 U482 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n437) );
  NOR2_X1 U483 ( .A1(n557), .A2(n423), .ZN(n582) );
  INV_X1 U484 ( .A(n576), .ZN(n360) );
  NAND2_X1 U485 ( .A1(n430), .A2(n429), .ZN(n359) );
  INV_X1 U486 ( .A(n644), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n431), .B(n524), .ZN(n430) );
  XOR2_X1 U488 ( .A(n459), .B(n458), .Z(n535) );
  XNOR2_X1 U489 ( .A(n414), .B(n410), .ZN(n465) );
  BUF_X1 U490 ( .A(n699), .Z(n708) );
  XNOR2_X1 U491 ( .A(n481), .B(n480), .ZN(n482) );
  NOR2_X1 U492 ( .A1(n602), .A2(n599), .ZN(n578) );
  NAND2_X1 U493 ( .A1(n370), .A2(n374), .ZN(n369) );
  AND2_X1 U494 ( .A1(n376), .A2(n372), .ZN(n371) );
  XNOR2_X1 U495 ( .A(n531), .B(n530), .ZN(n741) );
  XNOR2_X1 U496 ( .A(KEYINPUT32), .B(KEYINPUT65), .ZN(n530) );
  XNOR2_X1 U497 ( .A(n592), .B(n406), .ZN(n739) );
  INV_X1 U498 ( .A(KEYINPUT105), .ZN(n406) );
  INV_X1 U499 ( .A(n593), .ZN(n625) );
  INV_X1 U500 ( .A(n359), .ZN(n622) );
  NOR2_X1 U501 ( .A1(n610), .A2(n712), .ZN(n613) );
  NOR2_X1 U502 ( .A1(n703), .A2(n712), .ZN(n363) );
  NOR2_X1 U503 ( .A1(n712), .A2(n692), .ZN(n693) );
  XNOR2_X1 U504 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U505 ( .A(KEYINPUT6), .B(n555), .ZN(n525) );
  XNOR2_X1 U506 ( .A(G119), .B(KEYINPUT3), .ZN(n353) );
  XOR2_X1 U507 ( .A(G131), .B(G134), .Z(n354) );
  AND2_X1 U508 ( .A1(G210), .A2(n511), .ZN(n355) );
  AND2_X1 U509 ( .A1(n538), .A2(n519), .ZN(n356) );
  OR2_X1 U510 ( .A1(n368), .A2(G902), .ZN(n357) );
  XOR2_X1 U511 ( .A(KEYINPUT48), .B(KEYINPUT69), .Z(n358) );
  INV_X1 U512 ( .A(KEYINPUT44), .ZN(n392) );
  XNOR2_X2 U513 ( .A(n523), .B(KEYINPUT22), .ZN(n527) );
  NAND2_X1 U514 ( .A1(n359), .A2(n390), .ZN(n381) );
  INV_X1 U515 ( .A(n565), .ZN(n555) );
  AND2_X1 U516 ( .A1(n565), .A2(n360), .ZN(n556) );
  XNOR2_X1 U517 ( .A(n596), .B(n358), .ZN(n388) );
  NAND2_X1 U518 ( .A1(n388), .A2(n386), .ZN(n732) );
  XNOR2_X1 U519 ( .A(n363), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U520 ( .A1(n694), .A2(n368), .ZN(n364) );
  NAND2_X1 U521 ( .A1(n666), .A2(n356), .ZN(n376) );
  INV_X1 U522 ( .A(n666), .ZN(n370) );
  AND2_X1 U523 ( .A1(n373), .A2(n520), .ZN(n372) );
  NAND2_X1 U524 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U525 ( .A1(n378), .A2(n377), .ZN(n382) );
  NAND2_X1 U526 ( .A1(n545), .A2(n392), .ZN(n377) );
  NAND2_X1 U527 ( .A1(n379), .A2(n532), .ZN(n378) );
  NOR2_X1 U528 ( .A1(n381), .A2(n380), .ZN(n379) );
  INV_X1 U529 ( .A(n545), .ZN(n380) );
  NOR2_X2 U530 ( .A1(n716), .A2(n732), .ZN(n673) );
  XNOR2_X2 U531 ( .A(n389), .B(n546), .ZN(n716) );
  INV_X1 U532 ( .A(n581), .ZN(n393) );
  NAND2_X1 U533 ( .A1(n400), .A2(n538), .ZN(n523) );
  NAND2_X1 U534 ( .A1(n517), .A2(n399), .ZN(n397) );
  NAND2_X1 U535 ( .A1(n581), .A2(n399), .ZN(n398) );
  INV_X1 U536 ( .A(KEYINPUT0), .ZN(n399) );
  NAND2_X1 U537 ( .A1(n636), .A2(n408), .ZN(n407) );
  NAND2_X1 U538 ( .A1(n580), .A2(n600), .ZN(n636) );
  INV_X1 U539 ( .A(n553), .ZN(n644) );
  NAND2_X1 U540 ( .A1(n417), .A2(n582), .ZN(n563) );
  NAND2_X1 U541 ( .A1(n417), .A2(n351), .ZN(n682) );
  NAND2_X1 U542 ( .A1(n655), .A2(n417), .ZN(n669) );
  INV_X1 U543 ( .A(n558), .ZN(n602) );
  NAND2_X1 U544 ( .A1(n425), .A2(n424), .ZN(n426) );
  NOR2_X1 U545 ( .A1(n527), .A2(n600), .ZN(n542) );
  XNOR2_X1 U546 ( .A(KEYINPUT46), .B(KEYINPUT86), .ZN(n433) );
  XNOR2_X1 U547 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n434) );
  INV_X1 U548 ( .A(KEYINPUT90), .ZN(n478) );
  XNOR2_X1 U549 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U550 ( .A(KEYINPUT106), .ZN(n560) );
  XNOR2_X1 U551 ( .A(n503), .B(n497), .ZN(n498) );
  XNOR2_X1 U552 ( .A(n460), .B(n440), .ZN(n441) );
  XNOR2_X1 U553 ( .A(G475), .B(KEYINPUT13), .ZN(n443) );
  XNOR2_X1 U554 ( .A(n694), .B(n695), .ZN(n696) );
  XNOR2_X1 U555 ( .A(KEYINPUT101), .B(n574), .ZN(n628) );
  XNOR2_X1 U556 ( .A(n611), .B(KEYINPUT108), .ZN(n612) );
  XNOR2_X1 U557 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U558 ( .A(n435), .B(n502), .ZN(n439) );
  XNOR2_X1 U559 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U560 ( .A(n439), .B(n438), .Z(n442) );
  NOR2_X1 U561 ( .A1(G953), .A2(G237), .ZN(n496) );
  NAND2_X1 U562 ( .A1(G214), .A2(n496), .ZN(n440) );
  NOR2_X1 U563 ( .A1(G902), .A2(n700), .ZN(n444) );
  XNOR2_X1 U564 ( .A(G478), .B(KEYINPUT98), .ZN(n445) );
  XNOR2_X1 U565 ( .A(n445), .B(KEYINPUT99), .ZN(n459) );
  XNOR2_X1 U566 ( .A(n475), .B(KEYINPUT9), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U568 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n450) );
  XNOR2_X1 U569 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U570 ( .A(n452), .B(n451), .Z(n455) );
  NAND2_X1 U571 ( .A1(G234), .A2(n734), .ZN(n453) );
  XOR2_X1 U572 ( .A(KEYINPUT8), .B(n453), .Z(n463) );
  NAND2_X1 U573 ( .A1(G217), .A2(n463), .ZN(n454) );
  XNOR2_X1 U574 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U575 ( .A(n457), .B(n456), .ZN(n705) );
  INV_X1 U576 ( .A(n535), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n533), .A2(n522), .ZN(n591) );
  XNOR2_X1 U578 ( .A(n591), .B(KEYINPUT79), .ZN(n520) );
  XNOR2_X1 U579 ( .A(n460), .B(n476), .ZN(n725) );
  NAND2_X1 U580 ( .A1(G221), .A2(n463), .ZN(n464) );
  XNOR2_X1 U581 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U582 ( .A(n725), .B(n466), .ZN(n707) );
  NOR2_X1 U583 ( .A1(n707), .A2(G902), .ZN(n471) );
  XOR2_X1 U584 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n469) );
  NAND2_X1 U585 ( .A1(G234), .A2(n604), .ZN(n467) );
  XNOR2_X1 U586 ( .A(KEYINPUT20), .B(n467), .ZN(n472) );
  NAND2_X1 U587 ( .A1(n472), .A2(G217), .ZN(n468) );
  XNOR2_X1 U588 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U589 ( .A(n471), .B(n470), .ZN(n553) );
  NAND2_X1 U590 ( .A1(n472), .A2(G221), .ZN(n473) );
  XNOR2_X1 U591 ( .A(n473), .B(KEYINPUT21), .ZN(n552) );
  INV_X1 U592 ( .A(n552), .ZN(n643) );
  NAND2_X1 U593 ( .A1(G227), .A2(n734), .ZN(n479) );
  XNOR2_X1 U594 ( .A(n484), .B(KEYINPUT74), .ZN(n537) );
  XOR2_X1 U595 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n486) );
  XNOR2_X1 U596 ( .A(G137), .B(KEYINPUT93), .ZN(n485) );
  XNOR2_X1 U597 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U598 ( .A(KEYINPUT70), .ZN(n489) );
  NAND2_X1 U599 ( .A1(G101), .A2(n489), .ZN(n492) );
  NAND2_X1 U600 ( .A1(n490), .A2(KEYINPUT70), .ZN(n491) );
  AND2_X1 U601 ( .A1(n496), .A2(G210), .ZN(n497) );
  NOR2_X1 U602 ( .A1(n607), .A2(G902), .ZN(n499) );
  NAND2_X1 U603 ( .A1(n537), .A2(n525), .ZN(n501) );
  XOR2_X1 U604 ( .A(n504), .B(KEYINPUT16), .Z(n505) );
  NAND2_X1 U605 ( .A1(G224), .A2(n734), .ZN(n508) );
  NAND2_X1 U606 ( .A1(n687), .A2(n604), .ZN(n510) );
  NAND2_X1 U607 ( .A1(G214), .A2(n511), .ZN(n656) );
  NAND2_X1 U608 ( .A1(n558), .A2(n656), .ZN(n513) );
  INV_X1 U609 ( .A(KEYINPUT19), .ZN(n512) );
  NAND2_X1 U610 ( .A1(G234), .A2(G237), .ZN(n514) );
  XNOR2_X1 U611 ( .A(n514), .B(KEYINPUT14), .ZN(n515) );
  NAND2_X1 U612 ( .A1(G952), .A2(n515), .ZN(n672) );
  NOR2_X1 U613 ( .A1(G953), .A2(n672), .ZN(n551) );
  NAND2_X1 U614 ( .A1(G902), .A2(n515), .ZN(n547) );
  INV_X1 U615 ( .A(G898), .ZN(n715) );
  NAND2_X1 U616 ( .A1(G953), .A2(n715), .ZN(n719) );
  NOR2_X1 U617 ( .A1(n547), .A2(n719), .ZN(n516) );
  NOR2_X1 U618 ( .A1(n551), .A2(n516), .ZN(n517) );
  XOR2_X1 U619 ( .A(KEYINPUT34), .B(KEYINPUT80), .Z(n518) );
  XNOR2_X1 U620 ( .A(KEYINPUT72), .B(n518), .ZN(n519) );
  NOR2_X1 U621 ( .A1(n738), .A2(KEYINPUT67), .ZN(n532) );
  INV_X1 U622 ( .A(KEYINPUT66), .ZN(n524) );
  INV_X1 U623 ( .A(n352), .ZN(n600) );
  XOR2_X1 U624 ( .A(KEYINPUT81), .B(n525), .Z(n526) );
  NOR2_X1 U625 ( .A1(n644), .A2(n352), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT94), .ZN(n534) );
  NAND2_X1 U628 ( .A1(n534), .A2(n535), .ZN(n574) );
  NOR2_X1 U629 ( .A1(n535), .A2(n534), .ZN(n631) );
  INV_X1 U630 ( .A(n631), .ZN(n597) );
  NAND2_X1 U631 ( .A1(n574), .A2(n597), .ZN(n661) );
  XOR2_X1 U632 ( .A(n661), .B(KEYINPUT84), .Z(n584) );
  INV_X1 U633 ( .A(n555), .ZN(n647) );
  NAND2_X1 U634 ( .A1(n564), .A2(n538), .ZN(n536) );
  NOR2_X1 U635 ( .A1(n647), .A2(n536), .ZN(n619) );
  AND2_X1 U636 ( .A1(n537), .A2(n647), .ZN(n652) );
  NAND2_X1 U637 ( .A1(n538), .A2(n652), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n539), .B(KEYINPUT31), .ZN(n632) );
  NOR2_X1 U639 ( .A1(n619), .A2(n632), .ZN(n540) );
  NOR2_X1 U640 ( .A1(n584), .A2(n540), .ZN(n544) );
  NOR2_X1 U641 ( .A1(n525), .A2(n553), .ZN(n541) );
  NAND2_X1 U642 ( .A1(n542), .A2(n541), .ZN(n614) );
  INV_X1 U643 ( .A(n614), .ZN(n543) );
  XOR2_X1 U644 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n546) );
  NOR2_X1 U645 ( .A1(G900), .A2(n547), .ZN(n548) );
  NAND2_X1 U646 ( .A1(G953), .A2(n548), .ZN(n549) );
  XOR2_X1 U647 ( .A(KEYINPUT102), .B(n549), .Z(n550) );
  NOR2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n568) );
  NOR2_X1 U649 ( .A1(n568), .A2(n552), .ZN(n554) );
  NAND2_X1 U650 ( .A1(n554), .A2(n553), .ZN(n576) );
  XOR2_X1 U651 ( .A(KEYINPUT28), .B(n556), .Z(n557) );
  XNOR2_X1 U652 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n559) );
  NAND2_X1 U653 ( .A1(n662), .A2(n561), .ZN(n562) );
  XNOR2_X1 U654 ( .A(n563), .B(KEYINPUT42), .ZN(n743) );
  NAND2_X1 U655 ( .A1(n565), .A2(n656), .ZN(n566) );
  XNOR2_X1 U656 ( .A(n566), .B(KEYINPUT30), .ZN(n567) );
  NOR2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U658 ( .A1(n570), .A2(n569), .ZN(n588) );
  INV_X1 U659 ( .A(n657), .ZN(n571) );
  XNOR2_X1 U660 ( .A(n572), .B(KEYINPUT39), .ZN(n598) );
  XNOR2_X1 U661 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n579) );
  NAND2_X1 U662 ( .A1(n525), .A2(n628), .ZN(n575) );
  NOR2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n577), .A2(n656), .ZN(n599) );
  XOR2_X1 U665 ( .A(n579), .B(n578), .Z(n580) );
  XOR2_X1 U666 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n586) );
  NAND2_X1 U667 ( .A1(n393), .A2(n582), .ZN(n583) );
  XNOR2_X1 U668 ( .A(n583), .B(KEYINPUT82), .ZN(n593) );
  NOR2_X1 U669 ( .A1(n593), .A2(n584), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n602), .A2(n588), .ZN(n589) );
  XOR2_X1 U672 ( .A(KEYINPUT104), .B(n589), .Z(n590) );
  NOR2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n661), .A2(n625), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n594), .A2(KEYINPUT47), .ZN(n595) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n637) );
  OR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U678 ( .A(n601), .B(KEYINPUT43), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n639) );
  NOR2_X4 U680 ( .A1(n605), .A2(n604), .ZN(n699) );
  NAND2_X1 U681 ( .A1(n699), .A2(G472), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT107), .B(KEYINPUT62), .Z(n606) );
  XNOR2_X1 U683 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n609), .B(n608), .ZN(n610) );
  INV_X1 U685 ( .A(KEYINPUT63), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(G57) );
  XNOR2_X1 U687 ( .A(n614), .B(G101), .ZN(G3) );
  NAND2_X1 U688 ( .A1(n619), .A2(n628), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n615), .B(G104), .ZN(G6) );
  XOR2_X1 U690 ( .A(KEYINPUT27), .B(KEYINPUT110), .Z(n617) );
  XNOR2_X1 U691 ( .A(G107), .B(KEYINPUT26), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n617), .B(n616), .ZN(n618) );
  XOR2_X1 U693 ( .A(KEYINPUT109), .B(n618), .Z(n621) );
  NAND2_X1 U694 ( .A1(n619), .A2(n631), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(G9) );
  XOR2_X1 U696 ( .A(G110), .B(n622), .Z(G12) );
  XOR2_X1 U697 ( .A(G128), .B(KEYINPUT29), .Z(n624) );
  NAND2_X1 U698 ( .A1(n631), .A2(n625), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(G30) );
  NAND2_X1 U700 ( .A1(n625), .A2(n628), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT112), .ZN(n627) );
  XNOR2_X1 U702 ( .A(G146), .B(n627), .ZN(G48) );
  XOR2_X1 U703 ( .A(G113), .B(KEYINPUT113), .Z(n630) );
  NAND2_X1 U704 ( .A1(n632), .A2(n628), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(G15) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(KEYINPUT114), .ZN(n634) );
  XNOR2_X1 U708 ( .A(G116), .B(n634), .ZN(G18) );
  XOR2_X1 U709 ( .A(G125), .B(KEYINPUT37), .Z(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(G27) );
  XNOR2_X1 U711 ( .A(G134), .B(n637), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n638), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U713 ( .A(G140), .B(n639), .ZN(G42) );
  NAND2_X1 U714 ( .A1(n352), .A2(n640), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT50), .B(n642), .Z(n650) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U717 ( .A(KEYINPUT49), .B(n645), .Z(n646) );
  NOR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U719 ( .A(KEYINPUT116), .B(n648), .Z(n649) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U722 ( .A(n653), .B(KEYINPUT117), .Z(n654) );
  XNOR2_X1 U723 ( .A(KEYINPUT51), .B(n654), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U726 ( .A(KEYINPUT118), .B(n660), .Z(n664) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U729 ( .A(KEYINPUT119), .B(n665), .Z(n667) );
  NAND2_X1 U730 ( .A1(n667), .A2(n351), .ZN(n668) );
  NAND2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U732 ( .A(KEYINPUT52), .B(n670), .Z(n671) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n681) );
  XNOR2_X1 U734 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n676) );
  NAND2_X1 U735 ( .A1(n676), .A2(n732), .ZN(n675) );
  NAND2_X1 U736 ( .A1(KEYINPUT2), .A2(n673), .ZN(n674) );
  NAND2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U738 ( .A1(n676), .A2(n716), .ZN(n677) );
  XNOR2_X1 U739 ( .A(KEYINPUT85), .B(n677), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U743 ( .A1(G953), .A2(n684), .ZN(n686) );
  XNOR2_X1 U744 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n685) );
  XNOR2_X1 U745 ( .A(n686), .B(n685), .ZN(G75) );
  NAND2_X1 U746 ( .A1(n699), .A2(G210), .ZN(n691) );
  INV_X1 U747 ( .A(n687), .ZN(n689) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n688) );
  XNOR2_X1 U749 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U750 ( .A(KEYINPUT56), .B(n693), .ZN(G51) );
  NAND2_X1 U751 ( .A1(n708), .A2(G469), .ZN(n697) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n695) );
  NOR2_X1 U753 ( .A1(n712), .A2(n698), .ZN(G54) );
  NAND2_X1 U754 ( .A1(n699), .A2(G475), .ZN(n702) );
  XNOR2_X1 U755 ( .A(n700), .B(n434), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U757 ( .A1(G478), .A2(n708), .ZN(n704) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n712), .A2(n706), .ZN(G63) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT122), .ZN(n710) );
  NAND2_X1 U761 ( .A1(G217), .A2(n708), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(G66) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n713) );
  XOR2_X1 U765 ( .A(KEYINPUT61), .B(n713), .Z(n714) );
  NOR2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n718) );
  NOR2_X1 U767 ( .A1(G953), .A2(n716), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n724) );
  XOR2_X1 U769 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n722) );
  NAND2_X1 U770 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(G69) );
  XOR2_X1 U773 ( .A(n725), .B(KEYINPUT125), .Z(n726) );
  XNOR2_X1 U774 ( .A(n727), .B(n726), .ZN(n733) );
  XNOR2_X1 U775 ( .A(G227), .B(n733), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  XOR2_X1 U777 ( .A(KEYINPUT126), .B(n729), .Z(n730) );
  NOR2_X1 U778 ( .A1(n734), .A2(n730), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n731), .B(KEYINPUT127), .ZN(n737) );
  XNOR2_X1 U780 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U783 ( .A(G122), .B(n738), .Z(G24) );
  XNOR2_X1 U784 ( .A(G143), .B(n739), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n740), .B(KEYINPUT111), .ZN(G45) );
  XOR2_X1 U786 ( .A(n741), .B(G119), .Z(G21) );
  XNOR2_X1 U787 ( .A(G131), .B(n742), .ZN(G33) );
  XNOR2_X1 U788 ( .A(n743), .B(G137), .ZN(G39) );
endmodule

