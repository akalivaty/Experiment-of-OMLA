//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  AOI21_X1  g004(.A(G131), .B1(new_n189), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT64), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n190), .B(new_n193), .C1(G134), .C2(new_n192), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT0), .A3(G128), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT0), .B(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(new_n202), .A3(new_n207), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n196), .A2(new_n197), .B1(G131), .B2(new_n199), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n209), .B2(new_n206), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(new_n203), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n189), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n192), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n198), .A3(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n208), .A2(new_n210), .A3(new_n219), .ZN(new_n220));
  XOR2_X1   g034(.A(G116), .B(G119), .Z(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT2), .B(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT2), .B(G113), .Z(new_n224));
  XNOR2_X1  g038(.A(G116), .B(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT67), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n207), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n209), .B2(new_n206), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n231), .A3(new_n219), .ZN(new_n232));
  INV_X1    g046(.A(new_n227), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n220), .A2(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n235));
  OAI21_X1  g049(.A(new_n187), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n233), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n228), .A2(new_n208), .A3(new_n210), .A4(new_n219), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT70), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n219), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n209), .A2(new_n206), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n247), .B(KEYINPUT27), .Z(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n248), .B(new_n249), .Z(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n220), .A2(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n232), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n233), .A3(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n255), .A2(new_n238), .ZN(new_n256));
  INV_X1    g070(.A(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT29), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n244), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n220), .A2(new_n228), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n238), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n262), .B2(KEYINPUT28), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT29), .A3(new_n250), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(G472), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n255), .A2(new_n238), .A3(new_n250), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n272));
  NAND4_X1  g086(.A1(new_n255), .A2(new_n238), .A3(new_n250), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n244), .B1(new_n239), .B2(KEYINPUT70), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n187), .B(new_n235), .C1(new_n237), .C2(new_n238), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n257), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT71), .B(new_n257), .C1(new_n275), .C2(new_n276), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(G472), .A2(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n281), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  INV_X1    g099(.A(new_n274), .ZN(new_n286));
  INV_X1    g100(.A(new_n280), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT71), .B1(new_n245), .B2(new_n257), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n285), .B1(new_n289), .B2(new_n282), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n267), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G234), .ZN(new_n292));
  OAI21_X1  g106(.A(G217), .B1(new_n292), .B2(G902), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT72), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G137), .ZN(new_n296));
  INV_X1    g110(.A(G221), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n297), .A2(new_n292), .A3(G953), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n296), .B(new_n298), .Z(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G125), .B(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT16), .ZN(new_n302));
  INV_X1    g116(.A(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n304), .A2(KEYINPUT16), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(G146), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n302), .A2(KEYINPUT75), .A3(new_n305), .A4(G146), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n301), .A2(new_n212), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G128), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n312), .A2(G128), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(KEYINPUT23), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(G110), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  XNOR2_X1  g132(.A(G119), .B(G128), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n316), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n310), .A2(new_n311), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n305), .A4(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n302), .A2(new_n305), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n212), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n316), .A2(G110), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n318), .A2(new_n319), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n300), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n328), .A2(new_n331), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n321), .A3(new_n299), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n335), .A3(new_n265), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT25), .A4(new_n265), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n295), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n333), .ZN(new_n341));
  INV_X1    g155(.A(new_n335), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n294), .A2(G902), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n340), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G237), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G214), .ZN(new_n353));
  INV_X1    g167(.A(G143), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT90), .B1(new_n357), .B2(G131), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n359));
  INV_X1    g173(.A(G131), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n359), .B(new_n360), .C1(new_n355), .C2(new_n356), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n360), .A3(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n301), .A2(KEYINPUT19), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n301), .A2(KEYINPUT19), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n212), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n308), .A2(new_n309), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(KEYINPUT18), .A2(G131), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n304), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G146), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n311), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n355), .A2(new_n356), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT89), .A4(new_n377), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n364), .A2(new_n368), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT91), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  INV_X1    g201(.A(new_n385), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n308), .A2(new_n367), .A3(new_n309), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n362), .B2(new_n363), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n380), .A2(new_n381), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n387), .B(new_n388), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT17), .B1(new_n358), .B2(new_n361), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n328), .B(new_n393), .C1(new_n364), .C2(KEYINPUT17), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n380), .A2(new_n381), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n385), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n386), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(KEYINPUT92), .A3(new_n398), .A4(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n399), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT20), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n396), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n265), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G475), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT9), .B(G234), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(G217), .A3(new_n352), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G116), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n354), .A2(G128), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n211), .A2(G143), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n189), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT13), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n211), .A2(G143), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(KEYINPUT13), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(KEYINPUT93), .A3(new_n424), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n420), .B(new_n423), .C1(new_n430), .C2(new_n189), .ZN(new_n431));
  INV_X1    g245(.A(G116), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT14), .A3(G122), .ZN(new_n433));
  INV_X1    g247(.A(new_n418), .ZN(new_n434));
  OAI211_X1 g248(.A(G107), .B(new_n433), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g249(.A(new_n422), .ZN(new_n436));
  OAI21_X1  g250(.A(G134), .B1(new_n436), .B2(new_n427), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n437), .A2(new_n423), .B1(new_n419), .B2(new_n418), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n431), .A2(KEYINPUT94), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n430), .A2(new_n189), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n423), .A4(new_n420), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n417), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n442), .A3(new_n417), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n413), .B1(new_n446), .B2(new_n265), .ZN(new_n447));
  AOI211_X1 g261(.A(G902), .B(new_n412), .C1(new_n444), .C2(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(G234), .A2(G237), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G952), .A3(new_n352), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(G898), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(G902), .A3(G953), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT95), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n447), .A2(new_n448), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n406), .A2(new_n410), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n384), .A2(G107), .ZN(new_n463));
  AND2_X1   g277(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n464));
  NOR2_X1   g278(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n419), .B2(G104), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n419), .A2(G104), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT78), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n463), .B(new_n472), .C1(new_n465), .C2(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT79), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(KEYINPUT79), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(G101), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT80), .B(G101), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n471), .B2(new_n473), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT4), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n476), .A2(new_n482), .A3(G101), .A4(new_n477), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(KEYINPUT86), .A3(new_n233), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n384), .A2(G107), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n469), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n474), .B2(new_n479), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT87), .B(KEYINPUT5), .Z(new_n491));
  OR2_X1    g305(.A1(new_n221), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G113), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n432), .A2(G119), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n492), .A2(new_n495), .B1(new_n225), .B2(new_n224), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n471), .A2(KEYINPUT79), .A3(new_n473), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT79), .B1(new_n471), .B2(new_n473), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n499), .A2(new_n500), .A3(new_n487), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n227), .B1(new_n501), .B2(new_n482), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT86), .B1(new_n502), .B2(new_n484), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n462), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n484), .A2(new_n233), .A3(new_n485), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n507), .A2(new_n461), .A3(new_n497), .A4(new_n486), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(KEYINPUT6), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n206), .A2(G125), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(G125), .B2(new_n215), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT88), .B(G224), .Z(new_n512));
  OR2_X1    g326(.A1(new_n512), .A2(G953), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n511), .B(new_n513), .Z(new_n514));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n515), .B(new_n462), .C1(new_n498), .C2(new_n503), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(KEYINPUT7), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n511), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT5), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n495), .B1(new_n520), .B2(new_n221), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n226), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n490), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n461), .B(KEYINPUT8), .Z(new_n524));
  INV_X1    g338(.A(new_n490), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n496), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n519), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n508), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n460), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n517), .A2(new_n528), .A3(new_n460), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n458), .B(new_n459), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n297), .B1(new_n415), .B2(new_n265), .ZN(new_n533));
  INV_X1    g347(.A(G469), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n474), .A2(new_n479), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT4), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n207), .B(new_n485), .C1(new_n501), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n354), .A2(G146), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n213), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n214), .B(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n481), .A2(new_n540), .A3(new_n489), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT81), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT10), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n489), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n215), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(KEYINPUT81), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n537), .A2(new_n209), .A3(new_n543), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G140), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n352), .A2(G227), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT83), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT83), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n548), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n490), .A2(new_n215), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n201), .B1(new_n557), .B2(new_n541), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT12), .B(new_n201), .C1(new_n557), .C2(new_n541), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n554), .A2(KEYINPUT84), .A3(new_n556), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n537), .A2(new_n543), .A3(new_n547), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n201), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n548), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT85), .B1(new_n566), .B2(new_n551), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT85), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n568), .B(new_n552), .C1(new_n565), .C2(new_n548), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n563), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n553), .A2(KEYINPUT83), .B1(new_n561), .B2(new_n560), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT84), .B1(new_n571), .B2(new_n556), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n534), .B(new_n265), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n553), .B1(new_n201), .B2(new_n564), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n562), .A2(new_n548), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT82), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n562), .A2(KEYINPUT82), .A3(new_n548), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n574), .B1(new_n579), .B2(new_n551), .ZN(new_n580));
  OAI21_X1  g394(.A(G469), .B1(new_n580), .B2(G902), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n533), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n291), .A2(new_n350), .A3(new_n532), .A4(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n480), .ZN(G3));
  NAND2_X1  g398(.A1(new_n573), .A2(new_n581), .ZN(new_n585));
  INV_X1    g399(.A(new_n533), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G472), .B1(new_n281), .B2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n289), .A2(new_n282), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n350), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n459), .B(new_n455), .C1(new_n530), .C2(new_n529), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n446), .A2(new_n265), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n411), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n439), .A2(new_n442), .A3(new_n417), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n596), .B1(new_n597), .B2(new_n443), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n445), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n601), .A2(KEYINPUT33), .A3(new_n444), .A4(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(KEYINPUT96), .B(new_n596), .C1(new_n597), .C2(new_n443), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n411), .A2(G902), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n600), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n406), .A2(new_n410), .B1(new_n595), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n593), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n592), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT98), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT99), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT34), .B(G104), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n400), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n398), .B1(new_n397), .B2(new_n399), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n410), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n447), .A2(new_n448), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT100), .B1(new_n593), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n459), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n517), .A2(new_n528), .ZN(new_n623));
  INV_X1    g437(.A(new_n460), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n517), .A2(new_n528), .A3(new_n460), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n620), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n455), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n592), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  AND2_X1   g448(.A1(new_n588), .A2(new_n589), .ZN(new_n635));
  INV_X1    g449(.A(new_n340), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n334), .A2(new_n321), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n300), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n344), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n635), .A2(new_n532), .A3(new_n582), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(new_n641), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT32), .B1(new_n281), .B2(new_n283), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n289), .A2(new_n285), .A3(new_n282), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n645), .B1(new_n648), .B2(new_n267), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n582), .A2(new_n627), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n450), .B1(new_n453), .B2(G900), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n410), .B(new_n652), .C1(new_n616), .C2(new_n617), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n619), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT101), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NOR2_X1   g471(.A1(new_n256), .A2(new_n257), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n265), .B1(new_n262), .B2(new_n250), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n648), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n641), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n652), .B(KEYINPUT39), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n582), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n530), .A2(new_n529), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT38), .ZN(new_n669));
  INV_X1    g483(.A(new_n619), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n459), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n410), .B2(new_n406), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n668), .A2(KEYINPUT38), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n663), .A2(new_n666), .A3(new_n667), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  AND2_X1   g490(.A1(new_n608), .A2(new_n652), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n651), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  AOI21_X1  g493(.A(new_n591), .B1(new_n648), .B2(new_n267), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n265), .B1(new_n570), .B2(new_n572), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n534), .A2(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI221_X1 g497(.A(new_n265), .B1(KEYINPUT102), .B2(new_n534), .C1(new_n570), .C2(new_n572), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n586), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n680), .A2(new_n610), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND3_X1  g503(.A1(new_n631), .A2(new_n680), .A3(new_n686), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  AND4_X1   g505(.A1(new_n586), .A2(new_n627), .A3(new_n683), .A4(new_n684), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n649), .A2(new_n692), .A3(new_n458), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  OAI211_X1 g508(.A(new_n672), .B(new_n455), .C1(new_n529), .C2(new_n530), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n271), .B(new_n273), .C1(new_n263), .C2(new_n250), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n697), .A2(new_n698), .A3(new_n282), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n697), .B2(new_n282), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(KEYINPUT104), .B(G472), .C1(new_n281), .C2(G902), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n289), .A2(new_n265), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT104), .B1(new_n704), .B2(G472), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n346), .B(KEYINPUT105), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n696), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n692), .A3(new_n641), .A4(new_n677), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT106), .B(G125), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G27));
  NOR3_X1   g526(.A1(new_n530), .A2(new_n529), .A3(new_n622), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n585), .A2(new_n713), .A3(new_n586), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n680), .A2(new_n677), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n648), .A2(KEYINPUT108), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n646), .A2(new_n647), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n267), .A3(new_n720), .ZN(new_n721));
  AND4_X1   g535(.A1(KEYINPUT42), .A2(new_n582), .A3(new_n677), .A4(new_n713), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n707), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  NAND3_X1  g539(.A1(new_n680), .A2(new_n655), .A3(new_n714), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  XNOR2_X1  g541(.A(new_n713), .B(KEYINPUT112), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n607), .A2(new_n595), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n406), .A2(new_n410), .A3(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT43), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT43), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT111), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n590), .A2(new_n641), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT44), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n738), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n734), .A3(new_n741), .A4(new_n736), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n728), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n562), .A2(KEYINPUT82), .A3(new_n548), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT82), .B1(new_n562), .B2(new_n548), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n551), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n574), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(KEYINPUT45), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT110), .A4(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n580), .C2(KEYINPUT45), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n746), .B2(new_n747), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT109), .B1(new_n755), .B2(new_n534), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(G469), .A2(G902), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n573), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n586), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n743), .A2(new_n664), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n586), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n591), .A2(new_n677), .A3(new_n713), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n291), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND2_X1  g589(.A1(new_n721), .A2(new_n707), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n733), .A2(new_n450), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n586), .A2(new_n713), .A3(new_n684), .A4(new_n683), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(KEYINPUT121), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(KEYINPUT121), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n782), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n706), .A2(new_n777), .A3(new_n707), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n692), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n591), .A2(new_n450), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n662), .A2(new_n778), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n609), .ZN(new_n790));
  INV_X1    g604(.A(G952), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n791), .A3(G953), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n683), .A2(new_n684), .A3(new_n586), .A4(new_n622), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT118), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n795), .A2(KEYINPUT118), .B1(new_n673), .B2(new_n669), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n786), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n406), .A2(new_n410), .A3(new_n595), .A4(new_n607), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT104), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n588), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n641), .A3(new_n702), .A4(new_n701), .ZN(new_n806));
  OAI22_X1  g620(.A1(new_n789), .A2(new_n803), .B1(new_n779), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n786), .A2(new_n796), .A3(new_n797), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n794), .B1(new_n801), .B2(KEYINPUT120), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n586), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT47), .B1(new_n763), .B2(new_n586), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n683), .A2(new_n684), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n586), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n786), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n728), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n802), .B(new_n810), .C1(new_n815), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT51), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n817), .B1(new_n771), .B2(new_n814), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n802), .A4(new_n810), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n793), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n406), .A2(new_n410), .A3(new_n670), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n608), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n593), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n635), .A3(new_n350), .A4(new_n582), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n583), .A2(new_n829), .A3(new_n642), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n587), .A2(new_n531), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n590), .A2(new_n645), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n680), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n829), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n653), .A2(new_n670), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n714), .A2(new_n291), .A3(new_n641), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n726), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n723), .B2(new_n717), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n690), .A2(new_n708), .A3(new_n693), .A4(new_n687), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n582), .A2(new_n677), .A3(new_n713), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n806), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n806), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n837), .A2(new_n841), .A3(new_n843), .A4(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n649), .B(new_n650), .C1(new_n655), .C2(new_n677), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n672), .B(new_n652), .C1(new_n529), .C2(new_n530), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n661), .A2(new_n852), .A3(new_n582), .A4(new_n645), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n710), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n850), .A2(new_n710), .A3(new_n856), .A4(new_n853), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n825), .B1(new_n849), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n850), .A2(new_n710), .A3(new_n853), .A4(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n842), .B1(new_n836), .B2(new_n831), .ZN(new_n866));
  INV_X1    g680(.A(new_n840), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n724), .A2(new_n848), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n859), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n849), .A2(new_n825), .A3(new_n858), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n708), .A2(new_n693), .A3(new_n687), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n835), .A2(new_n583), .A3(new_n829), .A4(new_n642), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n835), .B1(new_n834), .B2(new_n829), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n690), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n724), .A2(new_n848), .A3(new_n867), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT116), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n868), .A2(new_n866), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n880), .A3(new_n865), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n872), .B1(new_n881), .B2(new_n825), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n824), .B(new_n871), .C1(new_n882), .C2(new_n870), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n791), .A2(new_n352), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n707), .A2(new_n586), .A3(new_n459), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n661), .A2(new_n730), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n673), .A2(new_n669), .B1(new_n813), .B2(KEYINPUT49), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n888), .C1(KEYINPUT49), .C2(new_n813), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT113), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(G75));
  NAND2_X1  g705(.A1(new_n859), .A2(new_n869), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n893), .A3(G210), .A4(G902), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n509), .A2(new_n516), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n514), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n265), .B1(new_n859), .B2(new_n869), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n901), .B2(G210), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n352), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n897), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n903), .A2(new_n907), .ZN(G51));
  XOR2_X1   g722(.A(new_n758), .B(KEYINPUT57), .Z(new_n909));
  AND3_X1   g723(.A1(new_n859), .A2(new_n869), .A3(new_n870), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n870), .B1(new_n859), .B2(new_n869), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n570), .A2(new_n572), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n901), .A2(new_n754), .A3(new_n752), .A4(new_n756), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n904), .B1(new_n914), .B2(new_n915), .ZN(G54));
  AND2_X1   g730(.A1(KEYINPUT58), .A2(G475), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n901), .A2(new_n397), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n397), .B1(new_n901), .B2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n904), .ZN(G60));
  NAND3_X1  g734(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n910), .B2(new_n911), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n905), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n871), .B1(new_n882), .B2(new_n870), .ZN(new_n927));
  INV_X1    g741(.A(new_n923), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(new_n921), .ZN(G63));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n859), .B2(new_n869), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n639), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n905), .B1(new_n934), .B2(new_n343), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n934), .A2(new_n343), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n905), .A4(new_n935), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n512), .B2(new_n451), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n866), .B2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n895), .B1(G898), .B2(new_n352), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  AND2_X1   g759(.A1(new_n850), .A2(new_n710), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n724), .A2(new_n946), .A3(new_n726), .ZN(new_n947));
  INV_X1    g761(.A(new_n672), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n776), .A2(new_n668), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n664), .B(new_n765), .C1(new_n743), .C2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n774), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n252), .A2(new_n254), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n365), .A2(new_n366), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(G900), .A2(G953), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n952), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n352), .B1(G227), .B2(G900), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n946), .A2(new_n961), .A3(new_n675), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT123), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n946), .B2(new_n675), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n771), .B2(new_n773), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n827), .A2(new_n622), .A3(new_n529), .A4(new_n530), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n680), .A2(new_n967), .A3(new_n582), .A4(new_n664), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT124), .Z(new_n969));
  NAND2_X1  g783(.A1(new_n766), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n958), .B(new_n960), .C1(new_n972), .C2(new_n955), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n766), .B2(new_n969), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n965), .B(new_n963), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n955), .B1(new_n977), .B2(new_n352), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n952), .A2(new_n956), .A3(new_n957), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n959), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n973), .A2(new_n980), .ZN(G72));
  INV_X1    g795(.A(new_n658), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n966), .A2(new_n971), .A3(new_n866), .ZN(new_n983));
  XOR2_X1   g797(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n951), .B2(new_n876), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n256), .A3(new_n257), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n905), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n982), .A2(new_n258), .A3(new_n986), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT127), .Z(new_n992));
  NOR2_X1   g806(.A1(new_n882), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n987), .A2(new_n990), .A3(new_n993), .ZN(G57));
endmodule


