

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800;

  OR2_X1 U369 ( .A1(n663), .A2(n425), .ZN(n424) );
  XNOR2_X1 U370 ( .A(G116), .B(G122), .ZN(n539) );
  XNOR2_X1 U371 ( .A(G110), .B(G107), .ZN(n366) );
  INV_X1 U372 ( .A(G125), .ZN(n507) );
  INV_X1 U373 ( .A(G128), .ZN(n486) );
  XNOR2_X1 U374 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n506) );
  XNOR2_X2 U375 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X2 U376 ( .A(n698), .B(n697), .ZN(n699) );
  AND2_X2 U377 ( .A1(n462), .A2(n357), .ZN(n461) );
  NAND2_X1 U378 ( .A1(n405), .A2(n408), .ZN(n365) );
  AND2_X2 U379 ( .A1(n406), .A2(n407), .ZN(n405) );
  INV_X1 U380 ( .A(KEYINPUT16), .ZN(n370) );
  XNOR2_X1 U381 ( .A(G143), .B(G113), .ZN(n549) );
  XNOR2_X1 U382 ( .A(G116), .B(G113), .ZN(n484) );
  XNOR2_X1 U383 ( .A(G101), .B(G104), .ZN(n526) );
  INV_X1 U384 ( .A(G902), .ZN(n426) );
  BUF_X1 U385 ( .A(G107), .Z(n445) );
  NAND2_X2 U386 ( .A1(n398), .A2(n397), .ZN(n626) );
  OR2_X1 U387 ( .A1(n603), .A2(n624), .ZN(n605) );
  OR2_X1 U388 ( .A1(n603), .A2(n741), .ZN(n393) );
  AND2_X2 U389 ( .A1(n443), .A2(n441), .ZN(n398) );
  NOR2_X2 U390 ( .A1(n374), .A2(n741), .ZN(n348) );
  INV_X4 U391 ( .A(G953), .ZN(n793) );
  XNOR2_X1 U392 ( .A(G110), .B(KEYINPUT23), .ZN(n468) );
  AND2_X2 U393 ( .A1(n421), .A2(n419), .ZN(n483) );
  AND2_X1 U394 ( .A1(n479), .A2(n358), .ZN(n475) );
  NAND2_X1 U395 ( .A1(n477), .A2(n476), .ZN(n474) );
  NAND2_X2 U396 ( .A1(n427), .A2(n424), .ZN(n603) );
  AND2_X1 U397 ( .A1(n478), .A2(n601), .ZN(n358) );
  XNOR2_X1 U398 ( .A(n417), .B(n504), .ZN(n510) );
  NOR2_X1 U399 ( .A1(n793), .A2(n590), .ZN(n591) );
  NAND2_X1 U400 ( .A1(G472), .A2(n426), .ZN(n425) );
  INV_X2 U401 ( .A(G104), .ZN(n485) );
  INV_X1 U402 ( .A(KEYINPUT31), .ZN(n349) );
  XNOR2_X1 U403 ( .A(KEYINPUT24), .B(G119), .ZN(n471) );
  NAND2_X1 U404 ( .A1(n383), .A2(n587), .ZN(n382) );
  AND2_X1 U405 ( .A1(n402), .A2(n399), .ZN(n379) );
  XNOR2_X1 U406 ( .A(n430), .B(KEYINPUT32), .ZN(n434) );
  XNOR2_X1 U407 ( .A(n570), .B(n569), .ZN(n579) );
  NOR2_X1 U408 ( .A1(n705), .A2(n536), .ZN(n403) );
  XNOR2_X1 U409 ( .A(n348), .B(KEYINPUT106), .ZN(n745) );
  XNOR2_X1 U410 ( .A(n393), .B(n453), .ZN(n392) );
  OR2_X1 U411 ( .A1(n374), .A2(n359), .ZN(n386) );
  AND2_X1 U412 ( .A1(n565), .A2(n566), .ZN(n719) );
  NAND2_X2 U413 ( .A1(n475), .A2(n474), .ZN(n516) );
  AND2_X1 U414 ( .A1(n413), .A2(n600), .ZN(n596) );
  AND2_X1 U415 ( .A1(n429), .A2(n428), .ZN(n427) );
  XNOR2_X1 U416 ( .A(n514), .B(n513), .ZN(n601) );
  XNOR2_X1 U417 ( .A(n501), .B(n500), .ZN(n511) );
  XNOR2_X1 U418 ( .A(n506), .B(n473), .ZN(n537) );
  XNOR2_X1 U419 ( .A(n485), .B(G122), .ZN(n544) );
  XNOR2_X1 U420 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n500) );
  XNOR2_X1 U421 ( .A(G125), .B(KEYINPUT17), .ZN(n459) );
  XNOR2_X2 U422 ( .A(G140), .B(KEYINPUT10), .ZN(n508) );
  XNOR2_X2 U423 ( .A(KEYINPUT4), .B(G146), .ZN(n518) );
  OR2_X2 U424 ( .A1(n351), .A2(n386), .ZN(n385) );
  XNOR2_X1 U425 ( .A(n391), .B(n452), .ZN(n351) );
  NAND2_X1 U426 ( .A1(n405), .A2(n408), .ZN(n694) );
  XNOR2_X1 U427 ( .A(n533), .B(n349), .ZN(n404) );
  BUF_X1 U428 ( .A(n440), .Z(n350) );
  XNOR2_X1 U429 ( .A(n391), .B(n452), .ZN(n611) );
  NAND2_X1 U430 ( .A1(n387), .A2(n385), .ZN(n352) );
  NAND2_X1 U431 ( .A1(n387), .A2(n385), .ZN(n396) );
  NAND2_X1 U432 ( .A1(n394), .A2(n392), .ZN(n391) );
  NOR2_X1 U433 ( .A1(n653), .A2(n646), .ZN(n647) );
  NAND2_X1 U434 ( .A1(n398), .A2(n397), .ZN(n353) );
  XNOR2_X1 U435 ( .A(n353), .B(KEYINPUT19), .ZN(n354) );
  XNOR2_X1 U436 ( .A(n626), .B(KEYINPUT19), .ZN(n615) );
  XNOR2_X1 U437 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X2 U438 ( .A(n522), .B(n369), .ZN(n775) );
  NAND2_X1 U439 ( .A1(n434), .A2(n433), .ZN(n581) );
  INV_X1 U440 ( .A(n672), .ZN(n433) );
  INV_X1 U441 ( .A(G237), .ZN(n491) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n545) );
  XOR2_X1 U443 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n503) );
  XNOR2_X1 U444 ( .A(n432), .B(KEYINPUT66), .ZN(n431) );
  NAND2_X1 U445 ( .A1(n581), .A2(KEYINPUT44), .ZN(n432) );
  NAND2_X1 U446 ( .A1(n447), .A2(KEYINPUT48), .ZN(n446) );
  AND2_X1 U447 ( .A1(n637), .A2(n442), .ZN(n439) );
  NAND2_X1 U448 ( .A1(n451), .A2(n719), .ZN(n627) );
  INV_X1 U449 ( .A(n624), .ZN(n451) );
  INV_X1 U450 ( .A(KEYINPUT30), .ZN(n453) );
  XNOR2_X1 U451 ( .A(n395), .B(n454), .ZN(n394) );
  INV_X1 U452 ( .A(KEYINPUT74), .ZN(n454) );
  XNOR2_X1 U453 ( .A(n471), .B(n470), .ZN(n469) );
  XNOR2_X1 U454 ( .A(n468), .B(n505), .ZN(n467) );
  INV_X1 U455 ( .A(G137), .ZN(n505) );
  NAND2_X1 U456 ( .A1(n793), .A2(G234), .ZN(n473) );
  NAND2_X1 U457 ( .A1(n537), .A2(G217), .ZN(n450) );
  XNOR2_X1 U458 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n547) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n548) );
  XNOR2_X1 U460 ( .A(n546), .B(n373), .ZN(n372) );
  INV_X1 U461 ( .A(KEYINPUT99), .ZN(n373) );
  XNOR2_X1 U462 ( .A(n415), .B(n438), .ZN(n414) );
  INV_X1 U463 ( .A(n518), .ZN(n438) );
  XNOR2_X1 U464 ( .A(n558), .B(n557), .ZN(n565) );
  INV_X1 U465 ( .A(KEYINPUT103), .ZN(n437) );
  INV_X1 U466 ( .A(n719), .ZN(n625) );
  INV_X1 U467 ( .A(KEYINPUT90), .ZN(n442) );
  OR2_X1 U468 ( .A1(n637), .A2(n442), .ZN(n441) );
  NAND2_X1 U469 ( .A1(n511), .A2(G217), .ZN(n417) );
  NAND2_X1 U470 ( .A1(n650), .A2(n649), .ZN(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT71), .B(G137), .ZN(n390) );
  NAND2_X1 U472 ( .A1(G237), .A2(G234), .ZN(n495) );
  INV_X1 U473 ( .A(KEYINPUT38), .ZN(n465) );
  NAND2_X1 U474 ( .A1(n510), .A2(n480), .ZN(n478) );
  NAND2_X1 U475 ( .A1(n524), .A2(G902), .ZN(n428) );
  XNOR2_X1 U476 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n520) );
  INV_X1 U477 ( .A(n627), .ZN(n638) );
  INV_X1 U478 ( .A(KEYINPUT73), .ZN(n452) );
  INV_X1 U479 ( .A(G469), .ZN(n455) );
  INV_X1 U480 ( .A(KEYINPUT0), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n663), .B(KEYINPUT62), .ZN(n664) );
  XNOR2_X1 U482 ( .A(n469), .B(n467), .ZN(n466) );
  XNOR2_X1 U483 ( .A(n449), .B(n448), .ZN(n657) );
  XNOR2_X1 U484 ( .A(n541), .B(n538), .ZN(n448) );
  XNOR2_X1 U485 ( .A(n372), .B(n544), .ZN(n554) );
  XNOR2_X1 U486 ( .A(n632), .B(KEYINPUT108), .ZN(n798) );
  NAND2_X1 U487 ( .A1(n579), .A2(n576), .ZN(n430) );
  AND2_X1 U488 ( .A1(n479), .A2(n478), .ZN(n355) );
  AND2_X1 U489 ( .A1(n413), .A2(n606), .ZN(n356) );
  AND2_X1 U490 ( .A1(n446), .A2(n797), .ZN(n357) );
  XNOR2_X1 U491 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n359) );
  XOR2_X1 U492 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n360) );
  BUF_X1 U493 ( .A(n755), .Z(n423) );
  AND2_X1 U494 ( .A1(KEYINPUT65), .A2(n761), .ZN(n361) );
  XNOR2_X1 U495 ( .A(n533), .B(KEYINPUT31), .ZN(n362) );
  XNOR2_X1 U496 ( .A(n459), .B(n458), .ZN(n457) );
  NAND2_X1 U497 ( .A1(n396), .A2(n719), .ZN(n599) );
  BUF_X1 U498 ( .A(n675), .Z(n422) );
  NAND2_X1 U499 ( .A1(n648), .A2(n760), .ZN(n363) );
  NAND2_X1 U500 ( .A1(n405), .A2(n408), .ZN(n364) );
  NOR2_X1 U501 ( .A1(n412), .A2(KEYINPUT65), .ZN(n410) );
  NAND2_X1 U502 ( .A1(n764), .A2(n411), .ZN(n412) );
  XNOR2_X1 U503 ( .A(n367), .B(n544), .ZN(n369) );
  XNOR2_X1 U504 ( .A(n525), .B(n370), .ZN(n367) );
  XNOR2_X2 U505 ( .A(n368), .B(n484), .ZN(n522) );
  XNOR2_X2 U506 ( .A(n371), .B(G119), .ZN(n368) );
  XNOR2_X2 U507 ( .A(G101), .B(KEYINPUT3), .ZN(n371) );
  NAND2_X1 U508 ( .A1(n379), .A2(n400), .ZN(n378) );
  XNOR2_X1 U509 ( .A(n378), .B(n437), .ZN(n377) );
  XNOR2_X1 U510 ( .A(n384), .B(n580), .ZN(n383) );
  NAND2_X1 U511 ( .A1(n374), .A2(n359), .ZN(n388) );
  NAND2_X1 U512 ( .A1(n374), .A2(n741), .ZN(n742) );
  XNOR2_X2 U513 ( .A(n612), .B(n465), .ZN(n374) );
  XNOR2_X2 U514 ( .A(n375), .B(n607), .ZN(n800) );
  NAND2_X1 U515 ( .A1(n740), .A2(n356), .ZN(n375) );
  XNOR2_X2 U516 ( .A(n376), .B(n360), .ZN(n740) );
  NAND2_X1 U517 ( .A1(n745), .A2(n743), .ZN(n376) );
  NAND2_X1 U518 ( .A1(n380), .A2(n377), .ZN(n436) );
  AND2_X1 U519 ( .A1(n381), .A2(n574), .ZN(n380) );
  NAND2_X1 U520 ( .A1(n675), .A2(KEYINPUT44), .ZN(n381) );
  XNOR2_X2 U521 ( .A(n481), .B(KEYINPUT35), .ZN(n675) );
  XNOR2_X2 U522 ( .A(n382), .B(KEYINPUT45), .ZN(n655) );
  NAND2_X1 U523 ( .A1(n435), .A2(n431), .ZN(n384) );
  AND2_X2 U524 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U525 ( .A1(n611), .A2(n359), .ZN(n389) );
  XNOR2_X1 U526 ( .A(n550), .B(n390), .ZN(n415) );
  XNOR2_X2 U527 ( .A(KEYINPUT70), .B(G131), .ZN(n550) );
  NAND2_X1 U528 ( .A1(n596), .A2(n595), .ZN(n395) );
  NAND2_X1 U529 ( .A1(n352), .A2(n722), .ZN(n670) );
  NAND2_X1 U530 ( .A1(n615), .A2(n499), .ZN(n444) );
  NAND2_X1 U531 ( .A1(n440), .A2(n439), .ZN(n397) );
  NAND2_X1 U532 ( .A1(n362), .A2(n536), .ZN(n399) );
  AND2_X1 U533 ( .A1(n401), .A2(n560), .ZN(n400) );
  NAND2_X1 U534 ( .A1(n705), .A2(n536), .ZN(n401) );
  NAND2_X1 U535 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U536 ( .A1(n363), .A2(n361), .ZN(n406) );
  NAND2_X1 U537 ( .A1(n412), .A2(KEYINPUT65), .ZN(n407) );
  NAND2_X1 U538 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U539 ( .A1(n363), .A2(n761), .ZN(n409) );
  NAND2_X1 U540 ( .A1(n769), .A2(n656), .ZN(n764) );
  AND2_X1 U541 ( .A1(n413), .A2(n731), .ZN(n534) );
  XNOR2_X1 U542 ( .A(n413), .B(KEYINPUT1), .ZN(n561) );
  XNOR2_X2 U543 ( .A(n456), .B(n455), .ZN(n413) );
  XNOR2_X2 U544 ( .A(n418), .B(n414), .ZN(n785) );
  XNOR2_X2 U545 ( .A(n517), .B(G134), .ZN(n418) );
  XNOR2_X2 U546 ( .A(n416), .B(n486), .ZN(n517) );
  XNOR2_X2 U547 ( .A(G143), .B(KEYINPUT76), .ZN(n416) );
  INV_X1 U548 ( .A(n601), .ZN(n725) );
  XNOR2_X1 U549 ( .A(n418), .B(n450), .ZN(n449) );
  NAND2_X1 U550 ( .A1(n532), .A2(n419), .ZN(n533) );
  NAND2_X1 U551 ( .A1(n419), .A2(n568), .ZN(n570) );
  AND2_X1 U552 ( .A1(n419), .A2(n535), .ZN(n705) );
  XNOR2_X2 U553 ( .A(n444), .B(n420), .ZN(n419) );
  INV_X1 U554 ( .A(n755), .ZN(n421) );
  XNOR2_X1 U555 ( .A(n472), .B(n466), .ZN(n509) );
  XNOR2_X1 U556 ( .A(n647), .B(KEYINPUT82), .ZN(n759) );
  NAND2_X1 U557 ( .A1(n663), .A2(n524), .ZN(n429) );
  XNOR2_X2 U558 ( .A(n785), .B(n523), .ZN(n663) );
  XNOR2_X2 U559 ( .A(n603), .B(KEYINPUT6), .ZN(n640) );
  INV_X1 U560 ( .A(n434), .ZN(n674) );
  XNOR2_X1 U561 ( .A(n436), .B(KEYINPUT87), .ZN(n435) );
  INV_X1 U562 ( .A(n597), .ZN(n440) );
  NAND2_X1 U563 ( .A1(n597), .A2(KEYINPUT90), .ZN(n443) );
  XNOR2_X1 U564 ( .A(n517), .B(n457), .ZN(n489) );
  OR2_X1 U565 ( .A1(n635), .A2(n636), .ZN(n460) );
  XNOR2_X2 U566 ( .A(n493), .B(n492), .ZN(n597) );
  NAND2_X1 U567 ( .A1(n633), .A2(n798), .ZN(n447) );
  INV_X1 U568 ( .A(n447), .ZN(n634) );
  NOR2_X2 U569 ( .A1(n689), .A2(G902), .ZN(n456) );
  XNOR2_X2 U570 ( .A(n785), .B(n530), .ZN(n689) );
  XNOR2_X2 U571 ( .A(KEYINPUT92), .B(KEYINPUT18), .ZN(n458) );
  AND2_X1 U572 ( .A1(n740), .A2(n748), .ZN(n756) );
  NAND2_X2 U573 ( .A1(n461), .A2(n460), .ZN(n464) );
  NAND2_X1 U574 ( .A1(n635), .A2(n463), .ZN(n462) );
  AND2_X1 U575 ( .A1(n634), .A2(n636), .ZN(n463) );
  XNOR2_X2 U576 ( .A(n464), .B(KEYINPUT84), .ZN(n653) );
  XNOR2_X2 U577 ( .A(G128), .B(KEYINPUT80), .ZN(n470) );
  NAND2_X1 U578 ( .A1(n537), .A2(G221), .ZN(n472) );
  NAND2_X1 U579 ( .A1(n676), .A2(n510), .ZN(n479) );
  NAND2_X1 U580 ( .A1(n355), .A2(n474), .ZN(n571) );
  NOR2_X1 U581 ( .A1(n510), .A2(n480), .ZN(n476) );
  INV_X1 U582 ( .A(n676), .ZN(n477) );
  INV_X1 U583 ( .A(n426), .ZN(n480) );
  NAND2_X1 U584 ( .A1(n482), .A2(n613), .ZN(n481) );
  XNOR2_X1 U585 ( .A(n483), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X2 U586 ( .A(n564), .B(n563), .ZN(n755) );
  XNOR2_X1 U587 ( .A(n659), .B(n658), .ZN(n661) );
  BUF_X1 U588 ( .A(n775), .Z(n777) );
  INV_X1 U589 ( .A(KEYINPUT63), .ZN(n667) );
  INV_X1 U590 ( .A(G110), .ZN(n671) );
  XNOR2_X2 U591 ( .A(G110), .B(G107), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n793), .A2(G224), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n518), .B(n487), .ZN(n488) );
  XNOR2_X1 U594 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U595 ( .A(n775), .B(n490), .ZN(n695) );
  XNOR2_X2 U596 ( .A(G902), .B(KEYINPUT15), .ZN(n649) );
  NAND2_X1 U597 ( .A1(n695), .A2(n649), .ZN(n493) );
  NAND2_X1 U598 ( .A1(n426), .A2(n491), .ZN(n494) );
  NAND2_X1 U599 ( .A1(n494), .A2(G210), .ZN(n492) );
  NAND2_X1 U600 ( .A1(n494), .A2(G214), .ZN(n637) );
  INV_X1 U601 ( .A(n637), .ZN(n741) );
  XOR2_X1 U602 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n496) );
  XNOR2_X1 U603 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U604 ( .A1(G952), .A2(n497), .ZN(n754) );
  OR2_X1 U605 ( .A1(n754), .A2(G953), .ZN(n594) );
  NAND2_X1 U606 ( .A1(G902), .A2(n497), .ZN(n590) );
  OR2_X1 U607 ( .A1(n793), .A2(G898), .ZN(n778) );
  OR2_X1 U608 ( .A1(n590), .A2(n778), .ZN(n498) );
  NAND2_X1 U609 ( .A1(n594), .A2(n498), .ZN(n499) );
  NAND2_X1 U610 ( .A1(n649), .A2(G234), .ZN(n501) );
  INV_X1 U611 ( .A(KEYINPUT75), .ZN(n502) );
  XNOR2_X1 U612 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U613 ( .A(n508), .B(n507), .ZN(n783) );
  XNOR2_X1 U614 ( .A(n783), .B(G146), .ZN(n555) );
  XNOR2_X1 U615 ( .A(n509), .B(n555), .ZN(n676) );
  NAND2_X1 U616 ( .A1(n511), .A2(G221), .ZN(n514) );
  INV_X1 U617 ( .A(KEYINPUT96), .ZN(n512) );
  XNOR2_X1 U618 ( .A(n512), .B(KEYINPUT21), .ZN(n513) );
  INV_X1 U619 ( .A(KEYINPUT68), .ZN(n515) );
  XNOR2_X2 U620 ( .A(n516), .B(n515), .ZN(n595) );
  BUF_X2 U621 ( .A(n595), .Z(n731) );
  NAND2_X1 U622 ( .A1(G210), .A2(n545), .ZN(n519) );
  XNOR2_X1 U623 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U624 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U625 ( .A(G472), .ZN(n524) );
  INV_X1 U626 ( .A(n603), .ZN(n728) );
  AND2_X1 U627 ( .A1(n731), .A2(n728), .ZN(n531) );
  XNOR2_X1 U628 ( .A(n366), .B(n526), .ZN(n529) );
  NAND2_X1 U629 ( .A1(n793), .A2(G227), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n527), .B(G140), .ZN(n528) );
  XNOR2_X1 U631 ( .A(n529), .B(n528), .ZN(n530) );
  BUF_X1 U632 ( .A(n561), .Z(n732) );
  NAND2_X1 U633 ( .A1(n531), .A2(n732), .ZN(n736) );
  INV_X1 U634 ( .A(n736), .ZN(n532) );
  AND2_X1 U635 ( .A1(n534), .A2(n603), .ZN(n535) );
  INV_X1 U636 ( .A(KEYINPUT98), .ZN(n536) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n538) );
  XOR2_X1 U638 ( .A(KEYINPUT102), .B(n445), .Z(n540) );
  XNOR2_X1 U639 ( .A(n540), .B(n539), .ZN(n541) );
  NAND2_X1 U640 ( .A1(n657), .A2(n426), .ZN(n543) );
  INV_X1 U641 ( .A(G478), .ZN(n542) );
  XNOR2_X1 U642 ( .A(n543), .B(n542), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n545), .A2(G214), .ZN(n546) );
  XNOR2_X1 U644 ( .A(n548), .B(n547), .ZN(n552) );
  XNOR2_X1 U645 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U646 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U647 ( .A(n554), .B(n553), .ZN(n556) );
  XNOR2_X1 U648 ( .A(n556), .B(n555), .ZN(n682) );
  NAND2_X1 U649 ( .A1(n682), .A2(n426), .ZN(n558) );
  XOR2_X1 U650 ( .A(KEYINPUT13), .B(G475), .Z(n557) );
  OR2_X1 U651 ( .A1(n566), .A2(n565), .ZN(n645) );
  NAND2_X1 U652 ( .A1(n625), .A2(n645), .ZN(n744) );
  INV_X1 U653 ( .A(KEYINPUT79), .ZN(n559) );
  XNOR2_X1 U654 ( .A(n744), .B(n559), .ZN(n560) );
  AND2_X1 U655 ( .A1(n731), .A2(n561), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n562), .A2(n640), .ZN(n564) );
  INV_X1 U657 ( .A(KEYINPUT33), .ZN(n563) );
  INV_X1 U658 ( .A(n565), .ZN(n567) );
  NOR2_X1 U659 ( .A1(n567), .A2(n566), .ZN(n613) );
  AND2_X1 U660 ( .A1(n567), .A2(n566), .ZN(n743) );
  AND2_X1 U661 ( .A1(n743), .A2(n601), .ZN(n568) );
  INV_X1 U662 ( .A(KEYINPUT22), .ZN(n569) );
  XNOR2_X1 U663 ( .A(n571), .B(KEYINPUT104), .ZN(n726) );
  OR2_X1 U664 ( .A1(n732), .A2(n726), .ZN(n572) );
  NOR2_X1 U665 ( .A1(n572), .A2(n640), .ZN(n573) );
  AND2_X1 U666 ( .A1(n579), .A2(n573), .ZN(n704) );
  INV_X1 U667 ( .A(n704), .ZN(n574) );
  NAND2_X1 U668 ( .A1(n732), .A2(n726), .ZN(n575) );
  NOR2_X1 U669 ( .A1(n575), .A2(n640), .ZN(n576) );
  NAND2_X1 U670 ( .A1(n603), .A2(n571), .ZN(n577) );
  NOR2_X1 U671 ( .A1(n732), .A2(n577), .ZN(n578) );
  AND2_X1 U672 ( .A1(n579), .A2(n578), .ZN(n672) );
  INV_X1 U673 ( .A(KEYINPUT86), .ZN(n580) );
  INV_X1 U674 ( .A(n581), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n582), .B(KEYINPUT88), .ZN(n586) );
  INV_X1 U676 ( .A(n422), .ZN(n584) );
  INV_X1 U677 ( .A(KEYINPUT44), .ZN(n583) );
  AND2_X1 U678 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U679 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U680 ( .A(n655), .B(KEYINPUT81), .ZN(n589) );
  INV_X1 U681 ( .A(n649), .ZN(n588) );
  NAND2_X1 U682 ( .A1(n589), .A2(n588), .ZN(n648) );
  INV_X1 U683 ( .A(G900), .ZN(n592) );
  NAND2_X1 U684 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U685 ( .A1(n594), .A2(n593), .ZN(n600) );
  BUF_X1 U686 ( .A(n597), .Z(n612) );
  INV_X1 U687 ( .A(KEYINPUT40), .ZN(n598) );
  XNOR2_X2 U688 ( .A(n599), .B(n598), .ZN(n673) );
  AND2_X1 U689 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U690 ( .A1(n571), .A2(n602), .ZN(n624) );
  INV_X1 U691 ( .A(KEYINPUT28), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n605), .B(n604), .ZN(n606) );
  INV_X1 U693 ( .A(KEYINPUT42), .ZN(n607) );
  NOR2_X2 U694 ( .A1(n673), .A2(n800), .ZN(n610) );
  XOR2_X1 U695 ( .A(KEYINPUT85), .B(KEYINPUT46), .Z(n608) );
  XNOR2_X1 U696 ( .A(n608), .B(KEYINPUT64), .ZN(n609) );
  XNOR2_X1 U697 ( .A(n610), .B(n609), .ZN(n635) );
  NAND2_X1 U698 ( .A1(n613), .A2(n350), .ZN(n614) );
  NOR2_X1 U699 ( .A1(n351), .A2(n614), .ZN(n714) );
  NAND2_X1 U700 ( .A1(n354), .A2(n356), .ZN(n710) );
  NOR2_X1 U701 ( .A1(n744), .A2(KEYINPUT79), .ZN(n616) );
  NOR2_X1 U702 ( .A1(n710), .A2(n616), .ZN(n617) );
  NOR2_X1 U703 ( .A1(n617), .A2(KEYINPUT47), .ZN(n622) );
  INV_X1 U704 ( .A(n744), .ZN(n619) );
  NOR2_X1 U705 ( .A1(KEYINPUT79), .A2(KEYINPUT47), .ZN(n618) );
  OR2_X1 U706 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U707 ( .A1(n710), .A2(n620), .ZN(n621) );
  NOR2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U709 ( .A1(n714), .A2(n623), .ZN(n633) );
  NOR2_X1 U710 ( .A1(n627), .A2(n353), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n628), .A2(n640), .ZN(n630) );
  XNOR2_X1 U712 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n631), .A2(n732), .ZN(n632) );
  INV_X1 U715 ( .A(KEYINPUT48), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U717 ( .A1(n639), .A2(n732), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n642), .B(KEYINPUT43), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n643), .A2(n612), .ZN(n644) );
  XOR2_X1 U721 ( .A(KEYINPUT105), .B(n644), .Z(n797) );
  INV_X1 U722 ( .A(n645), .ZN(n722) );
  INV_X1 U723 ( .A(n670), .ZN(n646) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n761) );
  NAND2_X1 U725 ( .A1(n759), .A2(KEYINPUT81), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n670), .A2(KEYINPUT2), .ZN(n651) );
  XOR2_X1 U727 ( .A(KEYINPUT77), .B(n651), .Z(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U729 ( .A(KEYINPUT83), .B(n654), .Z(n656) );
  BUF_X1 U730 ( .A(n655), .Z(n769) );
  NAND2_X1 U731 ( .A1(n365), .A2(G478), .ZN(n659) );
  INV_X1 U732 ( .A(n657), .ZN(n658) );
  INV_X1 U733 ( .A(G952), .ZN(n660) );
  AND2_X1 U734 ( .A1(n660), .A2(G953), .ZN(n701) );
  NOR2_X2 U735 ( .A1(n661), .A2(n701), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(KEYINPUT118), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n694), .A2(G472), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X2 U739 ( .A1(n666), .A2(n701), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(G57) );
  NAND2_X1 U741 ( .A1(n705), .A2(n719), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(G104), .ZN(G6) );
  XNOR2_X1 U743 ( .A(n670), .B(G134), .ZN(G36) );
  XNOR2_X1 U744 ( .A(n672), .B(n671), .ZN(G12) );
  XOR2_X1 U745 ( .A(n673), .B(G131), .Z(G33) );
  XOR2_X1 U746 ( .A(G119), .B(n674), .Z(G21) );
  XOR2_X1 U747 ( .A(n422), .B(G122), .Z(G24) );
  BUF_X1 U748 ( .A(n676), .Z(n677) );
  NAND2_X1 U749 ( .A1(n364), .A2(G217), .ZN(n678) );
  XNOR2_X1 U750 ( .A(n677), .B(n678), .ZN(n679) );
  NOR2_X1 U751 ( .A1(n679), .A2(n701), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n694), .A2(G475), .ZN(n684) );
  XNOR2_X1 U753 ( .A(KEYINPUT67), .B(KEYINPUT117), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n680), .B(KEYINPUT59), .ZN(n681) );
  XNOR2_X1 U755 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X2 U756 ( .A1(n685), .A2(n701), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U758 ( .A1(n364), .A2(G469), .ZN(n691) );
  XNOR2_X1 U759 ( .A(KEYINPUT115), .B(KEYINPUT57), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(KEYINPUT58), .ZN(n688) );
  XNOR2_X1 U761 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X2 U762 ( .A1(n692), .A2(n701), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT116), .ZN(G54) );
  NAND2_X1 U764 ( .A1(n365), .A2(G210), .ZN(n700) );
  BUF_X1 U765 ( .A(n695), .Z(n698) );
  XNOR2_X1 U766 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n696) );
  XOR2_X1 U767 ( .A(n696), .B(KEYINPUT55), .Z(n697) );
  XNOR2_X1 U768 ( .A(n700), .B(n699), .ZN(n702) );
  NOR2_X2 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U771 ( .A(G101), .B(n704), .Z(G3) );
  NAND2_X1 U772 ( .A1(n705), .A2(n722), .ZN(n707) );
  XOR2_X1 U773 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n706) );
  XNOR2_X1 U774 ( .A(n707), .B(n706), .ZN(n709) );
  XOR2_X1 U775 ( .A(n445), .B(KEYINPUT27), .Z(n708) );
  XNOR2_X1 U776 ( .A(n709), .B(n708), .ZN(G9) );
  XOR2_X1 U777 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n712) );
  INV_X1 U778 ( .A(n710), .ZN(n716) );
  NAND2_X1 U779 ( .A1(n716), .A2(n722), .ZN(n711) );
  XNOR2_X1 U780 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U781 ( .A(G128), .B(n713), .ZN(G30) );
  XNOR2_X1 U782 ( .A(G143), .B(n714), .ZN(n715) );
  XNOR2_X1 U783 ( .A(n715), .B(KEYINPUT111), .ZN(G45) );
  NAND2_X1 U784 ( .A1(n716), .A2(n719), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n717), .B(KEYINPUT112), .ZN(n718) );
  XNOR2_X1 U786 ( .A(G146), .B(n718), .ZN(G48) );
  XOR2_X1 U787 ( .A(G113), .B(KEYINPUT113), .Z(n721) );
  BUF_X1 U788 ( .A(n362), .Z(n723) );
  NAND2_X1 U789 ( .A1(n723), .A2(n719), .ZN(n720) );
  XNOR2_X1 U790 ( .A(n721), .B(n720), .ZN(G15) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U792 ( .A(n724), .B(G116), .ZN(G18) );
  NAND2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U794 ( .A(n727), .B(KEYINPUT49), .ZN(n729) );
  NOR2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U796 ( .A(n730), .B(KEYINPUT114), .ZN(n735) );
  NOR2_X1 U797 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U798 ( .A(KEYINPUT50), .B(n733), .Z(n734) );
  NAND2_X1 U799 ( .A1(n735), .A2(n734), .ZN(n737) );
  AND2_X1 U800 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U801 ( .A(KEYINPUT51), .B(n738), .ZN(n739) );
  NAND2_X1 U802 ( .A1(n740), .A2(n739), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U804 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U805 ( .A1(n747), .A2(n746), .ZN(n749) );
  INV_X1 U806 ( .A(n423), .ZN(n748) );
  NAND2_X1 U807 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U808 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U809 ( .A(KEYINPUT52), .B(n752), .Z(n753) );
  NOR2_X1 U810 ( .A1(n754), .A2(n753), .ZN(n757) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U812 ( .A1(n758), .A2(n793), .ZN(n767) );
  BUF_X1 U813 ( .A(n759), .Z(n760) );
  NAND2_X1 U814 ( .A1(n769), .A2(n760), .ZN(n762) );
  NAND2_X1 U815 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(KEYINPUT78), .ZN(n765) );
  AND2_X1 U817 ( .A1(n764), .A2(n765), .ZN(n766) );
  NOR2_X1 U818 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n768), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U820 ( .A1(n769), .A2(n793), .ZN(n774) );
  XOR2_X1 U821 ( .A(KEYINPUT61), .B(KEYINPUT119), .Z(n771) );
  NAND2_X1 U822 ( .A1(G224), .A2(G953), .ZN(n770) );
  XNOR2_X1 U823 ( .A(n771), .B(n770), .ZN(n772) );
  NAND2_X1 U824 ( .A1(n772), .A2(G898), .ZN(n773) );
  NAND2_X1 U825 ( .A1(n774), .A2(n773), .ZN(n781) );
  XNOR2_X1 U826 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n776) );
  XNOR2_X1 U827 ( .A(n777), .B(n776), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U829 ( .A(n781), .B(n780), .Z(n782) );
  XNOR2_X1 U830 ( .A(KEYINPUT122), .B(n782), .ZN(G69) );
  XOR2_X1 U831 ( .A(KEYINPUT123), .B(n783), .Z(n784) );
  XNOR2_X1 U832 ( .A(n785), .B(n784), .ZN(n791) );
  XNOR2_X1 U833 ( .A(n791), .B(G227), .ZN(n786) );
  XNOR2_X1 U834 ( .A(n786), .B(KEYINPUT125), .ZN(n787) );
  NAND2_X1 U835 ( .A1(n787), .A2(G900), .ZN(n788) );
  XOR2_X1 U836 ( .A(KEYINPUT126), .B(n788), .Z(n789) );
  NOR2_X1 U837 ( .A1(n793), .A2(n789), .ZN(n790) );
  XNOR2_X1 U838 ( .A(n790), .B(KEYINPUT127), .ZN(n796) );
  XNOR2_X1 U839 ( .A(n791), .B(KEYINPUT124), .ZN(n792) );
  XNOR2_X1 U840 ( .A(n760), .B(n792), .ZN(n794) );
  NAND2_X1 U841 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U842 ( .A1(n796), .A2(n795), .ZN(G72) );
  XNOR2_X1 U843 ( .A(G140), .B(n797), .ZN(G42) );
  XOR2_X1 U844 ( .A(G125), .B(n798), .Z(n799) );
  XNOR2_X1 U845 ( .A(KEYINPUT37), .B(n799), .ZN(G27) );
  XOR2_X1 U846 ( .A(n800), .B(G137), .Z(G39) );
endmodule

