//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  XOR2_X1   g000(.A(G110), .B(G122), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT81), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT72), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT72), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n194), .A3(new_n198), .A4(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(G101), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n191), .A2(new_n194), .A3(new_n203), .A4(new_n195), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT74), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n197), .A2(KEYINPUT73), .A3(G101), .A4(new_n199), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(KEYINPUT4), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G116), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT65), .B1(new_n208), .B2(G119), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n197), .A2(new_n217), .A3(G101), .A4(new_n199), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n207), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n195), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n190), .A2(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n204), .A2(KEYINPUT74), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n204), .A2(KEYINPUT74), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n214), .A2(new_n215), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n214), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n211), .A3(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G113), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n229), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n205), .A2(KEYINPUT75), .A3(new_n223), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n228), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n220), .A2(new_n238), .A3(KEYINPUT80), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT80), .B1(new_n220), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n189), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n220), .A2(new_n238), .A3(new_n188), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT6), .B(new_n189), .C1(new_n239), .C2(new_n240), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT0), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT0), .B(G128), .Z(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  OR2_X1    g066(.A1(KEYINPUT70), .A2(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT70), .A2(G125), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n247), .A2(new_n257), .A3(G128), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n259), .A3(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(G146), .C1(new_n249), .C2(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G224), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT82), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n266), .B(new_n269), .Z(new_n270));
  NAND2_X1  g084(.A1(new_n246), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT85), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n256), .A2(new_n265), .B1(new_n272), .B2(new_n269), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n236), .B1(new_n205), .B2(new_n223), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n235), .A2(KEYINPUT84), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n232), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n235), .A2(KEYINPUT84), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n231), .A2(KEYINPUT83), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n229), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n228), .A2(new_n237), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n276), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n187), .B(KEYINPUT8), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n275), .B(new_n244), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n271), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n271), .A2(new_n293), .A3(new_n291), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G214), .B1(G237), .B2(G902), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n298), .B(KEYINPUT79), .Z(new_n299));
  INV_X1    g113(.A(G221), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT9), .B(G234), .Z(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n289), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G137), .ZN(new_n306));
  INV_X1    g120(.A(G137), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT11), .A3(G134), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(G137), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G131), .ZN(new_n311));
  INV_X1    g125(.A(G131), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n306), .A2(new_n308), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(KEYINPUT64), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n315), .A3(G131), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n263), .B1(new_n228), .B2(new_n237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n205), .A2(new_n263), .A3(new_n223), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT12), .B(new_n318), .C1(new_n319), .C2(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n218), .A2(new_n252), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n207), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n264), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n228), .A2(new_n237), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n320), .A2(new_n329), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n331), .A3(new_n317), .A4(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n267), .A2(G227), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT77), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n326), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n318), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n333), .ZN(new_n345));
  INV_X1    g159(.A(new_n336), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI211_X1 g161(.A(KEYINPUT78), .B(new_n336), .C1(new_n344), .C2(new_n333), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n341), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G469), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n289), .ZN(new_n351));
  NAND2_X1  g165(.A1(G469), .A2(G902), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n326), .A2(new_n333), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n346), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n337), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n336), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n344), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(G469), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n297), .A2(new_n299), .A3(new_n303), .A4(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G143), .B1(new_n362), .B2(G214), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT17), .B(G131), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT90), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n368));
  INV_X1    g182(.A(G237), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n267), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n261), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n312), .B1(new_n371), .B2(new_n363), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n372), .B2(KEYINPUT17), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(KEYINPUT70), .A2(G125), .ZN(new_n375));
  NOR2_X1   g189(.A1(KEYINPUT70), .A2(G125), .ZN(new_n376));
  OAI21_X1  g190(.A(G140), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G125), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G140), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT16), .ZN(new_n382));
  INV_X1    g196(.A(G140), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n253), .A2(new_n382), .A3(new_n383), .A4(new_n254), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n259), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(G146), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT91), .B1(new_n374), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n371), .A2(new_n363), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n312), .ZN(new_n392));
  INV_X1    g206(.A(new_n372), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n366), .A2(KEYINPUT90), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n372), .A2(new_n368), .A3(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n387), .A4(new_n386), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n389), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT88), .B(G104), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n390), .B1(new_n406), .B2(new_n312), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n379), .B1(new_n255), .B2(G140), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n259), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n405), .A2(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n259), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT87), .B(new_n413), .C1(new_n408), .C2(new_n259), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n401), .A2(new_n404), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n404), .B1(new_n401), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n289), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G475), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n412), .A2(KEYINPUT19), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n408), .B2(KEYINPUT19), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n424), .A2(new_n259), .B1(new_n393), .B2(new_n392), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n425), .A2(new_n387), .B1(new_n411), .B2(new_n414), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n421), .B1(new_n426), .B2(new_n404), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n394), .B(new_n387), .C1(G146), .C2(new_n423), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n415), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n404), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(KEYINPUT89), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n416), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n432), .B2(new_n434), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n420), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT94), .ZN(new_n440));
  INV_X1    g254(.A(G478), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n301), .ZN(new_n444));
  INV_X1    g258(.A(G217), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n445), .A3(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  XNOR2_X1  g262(.A(G128), .B(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n305), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n208), .A2(G122), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n453), .A3(new_n193), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n193), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n249), .A2(G143), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n261), .A2(G128), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT13), .ZN(new_n459));
  OR3_X1    g273(.A1(new_n249), .A2(KEYINPUT13), .A3(G143), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n459), .A2(G134), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n448), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n452), .A2(G116), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n208), .A2(G122), .ZN(new_n464));
  OAI21_X1  g278(.A(G107), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n453), .A3(new_n193), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n465), .A2(new_n466), .B1(new_n305), .B2(new_n449), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n460), .A3(G134), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT92), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n449), .B(new_n305), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n193), .B1(new_n463), .B2(KEYINPUT14), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n451), .A2(new_n453), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(KEYINPUT14), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n466), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n471), .B1(new_n470), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n447), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n456), .A2(new_n461), .A3(new_n448), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT92), .B1(new_n467), .B2(new_n468), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT93), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n446), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n443), .B1(new_n486), .B2(new_n289), .ZN(new_n487));
  AOI211_X1 g301(.A(G902), .B(new_n442), .C1(new_n479), .C2(new_n485), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n440), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n477), .A2(new_n478), .A3(new_n447), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n446), .B1(new_n483), .B2(new_n484), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n289), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n442), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n289), .A3(new_n443), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(KEYINPUT94), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n439), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G952), .ZN(new_n498));
  AOI211_X1 g312(.A(G953), .B(new_n498), .C1(G234), .C2(G237), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT21), .B(G898), .Z(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n289), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT95), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n506));
  NOR4_X1   g320(.A1(new_n439), .A2(new_n496), .A3(new_n506), .A4(new_n503), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT96), .B1(new_n361), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n489), .A2(new_n495), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n432), .A2(new_n434), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n436), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(G475), .B2(new_n419), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n506), .B1(new_n515), .B2(new_n503), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n497), .A2(KEYINPUT95), .A3(new_n504), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n360), .A2(new_n303), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n293), .B1(new_n271), .B2(new_n291), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n294), .B(new_n290), .C1(new_n246), .C2(new_n270), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n299), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n518), .A2(new_n520), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n314), .A2(new_n252), .A3(new_n316), .ZN(new_n528));
  INV_X1    g342(.A(new_n216), .ZN(new_n529));
  INV_X1    g343(.A(new_n309), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n305), .A2(G137), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n263), .A2(new_n313), .A3(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n528), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n529), .B1(new_n528), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT28), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT67), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n534), .A2(KEYINPUT28), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(KEYINPUT28), .C1(new_n534), .C2(new_n535), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n362), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n533), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n528), .A2(KEYINPUT30), .A3(new_n533), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n216), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n528), .A2(new_n529), .A3(new_n533), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT66), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT66), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n558), .A3(KEYINPUT31), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(new_n556), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G472), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n289), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .A4(new_n289), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n541), .A2(new_n545), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n552), .A2(new_n546), .A3(new_n553), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT29), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n534), .A2(new_n535), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT68), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n553), .A2(KEYINPUT68), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(KEYINPUT28), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n572), .A2(KEYINPUT29), .A3(new_n545), .A4(new_n538), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n289), .ZN(new_n574));
  OAI21_X1  g388(.A(G472), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n564), .A2(new_n565), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n445), .B1(G234), .B2(new_n289), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n211), .A2(G128), .ZN(new_n579));
  NAND2_X1  g393(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n249), .A2(G119), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n581), .B(new_n583), .C1(KEYINPUT69), .C2(KEYINPUT23), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT71), .B(G110), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n582), .A2(new_n579), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT24), .B(G110), .Z(new_n587));
  OAI22_X1  g401(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n413), .A3(new_n387), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(G110), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n587), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n388), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT22), .B(G137), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n289), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n578), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n598), .A2(new_n599), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n605), .A2(G902), .A3(new_n577), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n576), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n509), .A2(new_n527), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT97), .B(G101), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G3));
  NAND2_X1  g426(.A1(new_n560), .A2(new_n289), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n614), .A2(new_n562), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n520), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n492), .A2(new_n441), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n486), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n479), .A2(new_n485), .A3(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n289), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(new_n441), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n439), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n298), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n295), .B2(new_n296), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n616), .A2(new_n504), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NOR2_X1   g445(.A1(new_n511), .A2(new_n436), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n420), .B1(new_n632), .B2(new_n438), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n510), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n616), .A2(new_n504), .A3(new_n626), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT100), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(G9));
  NAND2_X1  g452(.A1(new_n602), .A2(new_n603), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n577), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n593), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n577), .A2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n640), .A2(KEYINPUT101), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  INV_X1    g460(.A(new_n644), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n604), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n509), .A2(new_n527), .A3(new_n615), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  NAND4_X1  g466(.A1(new_n576), .A2(new_n303), .A3(new_n649), .A4(new_n360), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n298), .B1(new_n521), .B2(new_n522), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n502), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n499), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n633), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n510), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  AND2_X1   g478(.A1(new_n570), .A2(new_n571), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n289), .B1(new_n665), .B2(new_n545), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n552), .A2(new_n553), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n545), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n564), .A2(new_n565), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT102), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n523), .B(KEYINPUT38), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n659), .B(KEYINPUT39), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n520), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n510), .A2(new_n514), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n298), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n640), .A2(new_n644), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n674), .A2(new_n678), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  AND2_X1   g499(.A1(new_n576), .A2(new_n649), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n439), .A2(new_n622), .A3(new_n659), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n654), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n688), .A3(new_n689), .A4(new_n520), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n439), .A2(new_n622), .A3(new_n659), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n691), .B(new_n298), .C1(new_n521), .C2(new_n522), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT103), .B1(new_n653), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OAI211_X1 g509(.A(new_n504), .B(new_n298), .C1(new_n521), .C2(new_n522), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n608), .A2(new_n696), .A3(new_n623), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n349), .A2(new_n350), .A3(new_n289), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n350), .B1(new_n349), .B2(new_n289), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n698), .A2(new_n699), .A3(new_n302), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n701), .B(new_n703), .ZN(G15));
  NOR3_X1   g518(.A1(new_n604), .A2(new_n606), .A3(new_n503), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n626), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n576), .A2(new_n634), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n349), .A2(new_n289), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n303), .A3(new_n351), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n654), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n576), .A2(new_n634), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n705), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n686), .A3(new_n518), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n572), .A2(new_n720), .A3(new_n538), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n546), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n572), .B2(new_n538), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n557), .B(new_n555), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n561), .A3(new_n289), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n680), .A2(new_n614), .A3(new_n705), .A4(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n654), .A3(new_n711), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n452), .ZN(G24));
  NAND4_X1  g542(.A1(new_n691), .A2(new_n614), .A3(new_n682), .A4(new_n725), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n654), .A3(new_n711), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n378), .ZN(G27));
  NOR4_X1   g545(.A1(new_n608), .A2(new_n519), .A3(new_n297), .A4(new_n625), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT42), .B1(new_n732), .B2(new_n691), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n519), .A2(new_n297), .A3(new_n625), .ZN(new_n734));
  AND4_X1   g548(.A1(KEYINPUT42), .A2(new_n734), .A3(new_n609), .A4(new_n691), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n312), .ZN(G33));
  XNOR2_X1  g551(.A(new_n662), .B(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n732), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NOR2_X1   g554(.A1(new_n297), .A2(new_n625), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT43), .B1(new_n514), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n514), .A2(new_n622), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n615), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n682), .C1(new_n747), .C2(new_n746), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n742), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n354), .A2(KEYINPUT45), .A3(new_n358), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n354), .B2(new_n358), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n752), .B(G469), .C1(new_n756), .C2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n354), .A2(new_n358), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(G469), .A3(new_n753), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n352), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n351), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n303), .A3(new_n676), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n751), .B(new_n765), .C1(new_n750), .C2(new_n749), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n763), .B2(new_n303), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n742), .A2(new_n576), .A3(new_n607), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n762), .A2(new_n351), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT46), .B1(new_n761), .B2(new_n352), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n768), .B(new_n303), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n691), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NAND2_X1  g590(.A1(new_n498), .A2(new_n267), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n725), .A2(new_n614), .ZN(new_n778));
  INV_X1    g592(.A(new_n607), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n658), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n746), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n712), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(G952), .A3(new_n267), .ZN(new_n783));
  INV_X1    g597(.A(new_n672), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n741), .A2(new_n499), .A3(new_n700), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n783), .B1(new_n786), .B2(new_n624), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n746), .A2(new_n499), .A3(new_n700), .A4(new_n741), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n608), .B(new_n788), .C1(KEYINPUT117), .C2(KEYINPUT48), .ZN(new_n789));
  NOR2_X1   g603(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n698), .A2(new_n699), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n302), .ZN(new_n793));
  INV_X1    g607(.A(new_n774), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n769), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n741), .A3(new_n781), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT116), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n673), .A2(KEYINPUT113), .A3(new_n625), .A4(new_n700), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n523), .A2(KEYINPUT38), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n295), .A2(KEYINPUT38), .A3(new_n296), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n625), .B(new_n700), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n805), .A3(new_n781), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT115), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n811), .B2(new_n809), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n778), .A2(new_n682), .ZN(new_n813));
  INV_X1    g627(.A(new_n788), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n806), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n439), .A2(new_n622), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n786), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n796), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n799), .A2(new_n810), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n796), .B2(KEYINPUT116), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n815), .A2(new_n796), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n808), .A2(new_n809), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n787), .B(new_n791), .C1(new_n819), .C2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n799), .B1(new_n810), .B2(new_n818), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n820), .A3(new_n822), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT118), .A3(new_n787), .A4(new_n791), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n487), .A2(new_n488), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n623), .B1(new_n439), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n616), .A2(new_n504), .A3(new_n525), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n650), .A2(new_n610), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n727), .B1(new_n697), .B2(new_n700), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n716), .A2(new_n718), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n716), .A2(new_n836), .A3(KEYINPUT111), .A4(new_n718), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n734), .A2(new_n813), .A3(new_n691), .ZN(new_n842));
  INV_X1    g656(.A(new_n661), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n741), .A2(KEYINPUT112), .A3(new_n832), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n523), .A2(new_n832), .A3(new_n298), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n661), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n739), .B(new_n842), .C1(new_n653), .C2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n730), .B1(new_n655), .B2(new_n662), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n681), .A2(new_n523), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n682), .A2(new_n660), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n520), .A3(new_n671), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n694), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n850), .A2(new_n694), .A3(KEYINPUT52), .A4(new_n853), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n736), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n841), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n736), .B(new_n835), .C1(new_n839), .C2(new_n840), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n863), .B2(new_n858), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n835), .A2(new_n736), .A3(new_n837), .A4(new_n861), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n860), .A2(new_n861), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n777), .B1(new_n831), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT110), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n779), .A2(new_n745), .A3(new_n524), .A4(new_n302), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n784), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n792), .B(KEYINPUT49), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n873), .A2(new_n872), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n874), .A2(new_n673), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n871), .A2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n867), .A2(new_n289), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(G210), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n246), .B(new_n270), .Z(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n880), .B2(new_n881), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n267), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G51));
  NAND2_X1  g701(.A1(new_n352), .A2(KEYINPUT57), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n352), .A2(KEYINPUT57), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n867), .A2(new_n868), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n866), .A2(new_n858), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n864), .A2(new_n891), .A3(KEYINPUT54), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n349), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n879), .A2(G469), .A3(new_n756), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n886), .B1(new_n894), .B2(new_n895), .ZN(G54));
  INV_X1    g710(.A(new_n886), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  INV_X1    g712(.A(new_n432), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n860), .A2(new_n861), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n866), .A2(new_n858), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND4_X1   g718(.A1(KEYINPUT58), .A2(new_n904), .A3(G475), .A4(G902), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n905), .B2(new_n432), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n899), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n900), .B1(new_n906), .B2(new_n907), .ZN(G60));
  XNOR2_X1  g722(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n441), .A2(new_n289), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n909), .B(new_n910), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n870), .A2(new_n912), .B1(new_n620), .B2(new_n619), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n619), .A2(new_n620), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n914), .B(new_n911), .C1(new_n915), .C2(new_n869), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n913), .A2(new_n916), .A3(new_n886), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT123), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n919), .B(new_n920), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n605), .B1(new_n867), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n642), .B(new_n921), .C1(new_n864), .C2(new_n891), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n897), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n925), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT61), .B1(new_n925), .B2(KEYINPUT121), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(G66));
  INV_X1    g742(.A(new_n841), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n267), .B1(new_n500), .B2(G224), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n929), .A2(new_n267), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  INV_X1    g747(.A(new_n246), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(G898), .B2(new_n267), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  NAND2_X1  g750(.A1(new_n550), .A2(new_n551), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT125), .Z(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n424), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n766), .A2(new_n775), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n850), .A2(new_n694), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n765), .A2(new_n609), .A3(new_n851), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n940), .A2(new_n943), .A3(new_n859), .A4(new_n739), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n944), .B2(new_n267), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(G227), .B2(new_n267), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n732), .A2(new_n676), .A3(new_n833), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT62), .B1(new_n941), .B2(new_n684), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n941), .A2(KEYINPUT62), .A3(new_n684), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n940), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n267), .A3(new_n939), .ZN(new_n951));
  INV_X1    g765(.A(G227), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n656), .B1(new_n939), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n946), .B(new_n951), .C1(new_n267), .C2(new_n953), .ZN(G72));
  XNOR2_X1  g768(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n561), .A2(new_n289), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n950), .B2(new_n929), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n886), .B1(new_n958), .B2(new_n669), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n944), .B2(new_n929), .ZN(new_n960));
  INV_X1    g774(.A(new_n567), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n862), .A2(new_n864), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(new_n567), .A3(new_n668), .A4(new_n957), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n959), .A2(new_n962), .A3(new_n964), .ZN(G57));
endmodule


