//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT1), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n202), .B2(new_n203), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n207), .C1(new_n209), .C2(KEYINPUT66), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT67), .B(G113gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n204), .B(new_n208), .C1(new_n211), .C2(new_n203), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n217), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n225), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT28), .ZN(new_n228));
  AND4_X1   g027(.A1(new_n220), .A2(new_n222), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(new_n225), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n225), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n243), .B(new_n230), .C1(new_n231), .C2(new_n225), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n242), .A2(new_n233), .A3(new_n234), .A4(new_n244), .ZN(new_n245));
  AND4_X1   g044(.A1(KEYINPUT25), .A2(new_n236), .A3(new_n237), .A4(new_n239), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n240), .A2(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n214), .B1(new_n229), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n241), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n220), .A2(new_n222), .A3(new_n226), .A4(new_n228), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n213), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G227gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT34), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n254), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT32), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n257), .A3(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n248), .A2(new_n253), .A3(new_n266), .A4(new_n257), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT33), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  XOR2_X1   g068(.A(G15gat), .B(G43gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G71gat), .B(G99gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n260), .ZN(new_n275));
  AOI221_X4 g074(.A(new_n263), .B1(KEYINPUT33), .B2(new_n272), .C1(new_n265), .C2(new_n267), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n275), .ZN(new_n278));
  INV_X1    g077(.A(new_n268), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n265), .A2(new_n267), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT33), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n282), .A3(new_n272), .ZN(new_n283));
  INV_X1    g082(.A(new_n276), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n262), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n284), .A3(new_n278), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n261), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(KEYINPUT36), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT22), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n292), .A2(new_n293), .B1(G211gat), .B2(G218gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n292), .B2(new_n293), .ZN(new_n295));
  XNOR2_X1  g094(.A(G197gat), .B(G204gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G155gat), .B(G162gat), .Z(new_n301));
  XNOR2_X1  g100(.A(G141gat), .B(G148gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT75), .B(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G155gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT76), .B1(new_n305), .B2(KEYINPUT2), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n307), .B(new_n308), .C1(new_n304), .C2(G155gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n312));
  OR2_X1    g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n318), .A2(new_n319), .A3(new_n301), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n318), .B2(new_n301), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n310), .B(new_n311), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT79), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n301), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n319), .A3(new_n301), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n311), .A4(new_n310), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n300), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n310), .B1(new_n320), .B2(new_n321), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(KEYINPUT77), .A3(new_n310), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n311), .B1(new_n299), .B2(KEYINPUT29), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OR3_X1    g138(.A1(new_n332), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n338), .A2(new_n334), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n333), .B1(new_n332), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT31), .B(G50gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G22gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(KEYINPUT81), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n350), .B2(new_n346), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n351), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n340), .A2(new_n342), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n213), .B(KEYINPUT78), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n323), .B2(new_n329), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n327), .A2(new_n310), .A3(new_n214), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT80), .B1(new_n360), .B2(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(new_n334), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n214), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n361), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n359), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT5), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n213), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n336), .A2(new_n337), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n360), .ZN(new_n374));
  INV_X1    g173(.A(new_n368), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n364), .A3(new_n214), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n357), .A2(new_n358), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT0), .ZN(new_n384));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n386), .A3(new_n381), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n386), .B1(new_n377), .B2(new_n381), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G226gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n256), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n251), .A2(new_n252), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n331), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n395), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n300), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n299), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n406), .A2(KEYINPUT71), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(KEYINPUT71), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n406), .A2(new_n408), .ZN(new_n411));
  INV_X1    g210(.A(new_n405), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n402), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n355), .B1(new_n393), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT36), .B1(new_n286), .B2(new_n289), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n291), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n374), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n368), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(KEYINPUT39), .C1(new_n379), .C2(new_n368), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n386), .B(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n378), .A2(new_n366), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n359), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT39), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n375), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT40), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n423), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n382), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n422), .A2(KEYINPUT40), .A3(new_n423), .A4(new_n427), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n430), .A2(new_n415), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n369), .A2(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n423), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n388), .B1(new_n391), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n400), .A2(new_n402), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n412), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n409), .B(new_n407), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n434), .B(new_n355), .C1(new_n437), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT6), .B1(new_n435), .B2(new_n386), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n448), .A2(new_n432), .B1(KEYINPUT6), .B2(new_n392), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n415), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n437), .A2(KEYINPUT83), .A3(new_n416), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n352), .A2(new_n354), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n286), .B2(new_n289), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n289), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n261), .B1(new_n287), .B2(new_n288), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n355), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n393), .A2(new_n416), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT35), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n419), .A2(new_n446), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462));
  INV_X1    g261(.A(G8gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT16), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(G1gat), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n466), .B2(KEYINPUT88), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(G1gat), .B2(new_n464), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G50gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G43gat), .ZN(new_n471));
  INV_X1    g270(.A(G43gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G50gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT15), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n475));
  INV_X1    g274(.A(G29gat), .ZN(new_n476));
  INV_X1    g275(.A(G36gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n480), .A2(new_n481), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(KEYINPUT84), .A3(new_n479), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n472), .A2(G50gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n470), .A2(G43gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G29gat), .A2(G36gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n474), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n479), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n492));
  NOR2_X1   g291(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n477), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT17), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n484), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n484), .B2(new_n497), .ZN(new_n501));
  NOR3_X1   g300(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n481), .B1(new_n491), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n483), .A3(new_n489), .ZN(new_n504));
  INV_X1    g303(.A(new_n474), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n495), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n494), .B1(new_n493), .B2(new_n477), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n479), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n474), .A2(new_n489), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n488), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT86), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n501), .A2(new_n498), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n501), .A2(KEYINPUT87), .A3(new_n512), .A4(new_n498), .ZN(new_n516));
  AOI211_X1 g315(.A(new_n469), .B(new_n499), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n501), .A2(new_n512), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(new_n469), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT18), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n462), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n516), .ZN(new_n524));
  INV_X1    g323(.A(new_n469), .ZN(new_n525));
  INV_X1    g324(.A(new_n499), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  AOI211_X1 g327(.A(new_n528), .B(new_n519), .C1(new_n520), .C2(new_n469), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT89), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n518), .B(KEYINPUT13), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n520), .A2(new_n469), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n520), .A2(new_n469), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n527), .A2(new_n521), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n528), .ZN(new_n538));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G197gat), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT11), .B(G169gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT12), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n531), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n531), .B2(new_n538), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n461), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G85gat), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT93), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT7), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n553), .B(new_n556), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n562), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n557), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n553), .B1(new_n570), .B2(new_n556), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n524), .A2(new_n526), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT92), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT41), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(new_n520), .B2(new_n572), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(KEYINPUT95), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n576), .A2(new_n577), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n581), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n579), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n584), .A2(new_n585), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(KEYINPUT94), .A3(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n574), .A2(new_n594), .A3(new_n579), .A4(new_n590), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n599));
  AND2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(KEYINPUT9), .ZN(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(G71gat), .A2(G78gat), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n604), .A2(KEYINPUT90), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G57gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G64gat), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G57gat), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n604), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  AOI21_X1  g421(.A(new_n469), .B1(KEYINPUT21), .B2(new_n614), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n622), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n565), .A2(KEYINPUT96), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n614), .B(new_n630), .C1(new_n566), .C2(new_n571), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n556), .B1(new_n563), .B2(new_n564), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n552), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n605), .A2(new_n613), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n565), .B(new_n633), .C1(new_n634), .C2(KEYINPUT96), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT10), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n631), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n628), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n638), .A2(new_n640), .A3(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n598), .A2(new_n626), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n548), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n393), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g451(.A1(new_n650), .A2(new_n416), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT98), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G8gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n463), .B2(new_n653), .ZN(new_n657));
  MUX2_X1   g456(.A(new_n656), .B(new_n657), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g457(.A1(new_n286), .A2(new_n289), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT36), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n290), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n650), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n659), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n650), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n355), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n591), .A2(new_n589), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n583), .B2(new_n582), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n673), .A2(new_n585), .B1(new_n593), .B2(new_n596), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n461), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n455), .A2(new_n460), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n459), .A2(new_n453), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n446), .A2(new_n677), .A3(new_n290), .A4(new_n661), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n598), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n648), .B(KEYINPUT101), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n625), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n622), .B(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n683), .A2(new_n547), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n393), .ZN(new_n688));
  INV_X1    g487(.A(new_n648), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n598), .A2(new_n626), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT99), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n548), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n393), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n476), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n692), .A2(KEYINPUT100), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT100), .B1(new_n692), .B2(new_n694), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n688), .B1(new_n698), .B2(new_n699), .ZN(G1328gat));
  NOR3_X1   g499(.A1(new_n692), .A2(G36gat), .A3(new_n416), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  OAI21_X1  g501(.A(G36gat), .B1(new_n687), .B2(new_n416), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1329gat));
  NAND4_X1  g503(.A1(new_n675), .A2(new_n662), .A3(new_n680), .A4(new_n686), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G43gat), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT47), .B1(new_n706), .B2(KEYINPUT102), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n659), .A2(new_n472), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n692), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n707), .B(new_n709), .ZN(G1330gat));
  NAND4_X1  g509(.A1(new_n675), .A2(new_n453), .A3(new_n680), .A4(new_n686), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n548), .A2(new_n470), .A3(new_n453), .A4(new_n691), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT48), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n714), .B(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n546), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n531), .A2(new_n538), .A3(new_n544), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n598), .A3(new_n626), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n683), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT104), .B1(new_n461), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n679), .A2(new_n724), .A3(new_n683), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n393), .B(KEYINPUT105), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n608), .ZN(G1332gat));
  INV_X1    g528(.A(new_n726), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n415), .B1(new_n731), .B2(new_n610), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT106), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n610), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n723), .A2(new_n725), .A3(new_n659), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT107), .ZN(new_n738));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n725), .A3(new_n740), .A4(new_n659), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(G71gat), .A3(new_n662), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT50), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n453), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g549(.A(KEYINPUT108), .B1(new_n720), .B2(new_n685), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n547), .A2(new_n626), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n689), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n675), .A2(new_n693), .A3(new_n680), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G85gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n674), .B1(new_n676), .B2(new_n678), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n674), .B(new_n755), .C1(new_n676), .C2(new_n678), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(KEYINPUT51), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT109), .B1(new_n761), .B2(KEYINPUT51), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n693), .A2(new_n554), .A3(new_n648), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n758), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT110), .B(new_n758), .C1(new_n764), .C2(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1336gat));
  NAND4_X1  g569(.A1(new_n675), .A2(new_n415), .A3(new_n680), .A4(new_n756), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n761), .B2(KEYINPUT111), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n754), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT51), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n416), .A2(new_n682), .A3(G92gat), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n762), .B2(new_n763), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(new_n771), .B2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n681), .A2(new_n662), .A3(new_n756), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G99gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n689), .A2(G99gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n659), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n764), .B2(new_n790), .ZN(G1338gat));
  NAND4_X1  g590(.A1(new_n675), .A2(new_n453), .A3(new_n680), .A4(new_n756), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT53), .B1(new_n792), .B2(G106gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n355), .A2(new_n682), .A3(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n764), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n792), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n774), .A2(new_n777), .A3(new_n794), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT113), .B1(new_n792), .B2(G106gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(G1339gat));
  AOI21_X1  g601(.A(new_n518), .B1(new_n527), .B2(new_n535), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n534), .A2(new_n535), .A3(new_n533), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n542), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n719), .A2(new_n648), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(new_n629), .C1(new_n636), .C2(new_n637), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n645), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n628), .B(new_n810), .C1(new_n639), .C2(KEYINPUT10), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n638), .A3(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n647), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT55), .B1(new_n809), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT114), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n809), .A2(new_n812), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n647), .A4(new_n813), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n806), .B1(new_n547), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n674), .ZN(new_n824));
  INV_X1    g623(.A(new_n822), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n825), .A2(new_n719), .A3(new_n598), .A4(new_n805), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n626), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n721), .A2(new_n689), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n453), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(new_n693), .A3(new_n416), .A4(new_n659), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n547), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n727), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n454), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT115), .B1(new_n833), .B2(new_n454), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n416), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n720), .A2(new_n211), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n831), .B2(new_n682), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n648), .A2(new_n203), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT116), .Z(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n836), .B2(new_n841), .ZN(G1341gat));
  NOR2_X1   g641(.A1(new_n626), .A2(G127gat), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n416), .B(new_n843), .C1(new_n834), .C2(new_n835), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n831), .A2(new_n626), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n206), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n844), .B(new_n848), .C1(new_n206), .C2(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1342gat));
  NOR3_X1   g649(.A1(new_n674), .A2(G134gat), .A3(new_n415), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n834), .B2(new_n835), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n831), .B2(new_n674), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  NOR3_X1   g655(.A1(new_n662), .A2(new_n415), .A3(new_n355), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n833), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(G141gat), .A3(new_n547), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n828), .A2(new_n829), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n453), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n720), .A2(new_n598), .A3(new_n626), .A4(new_n648), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n719), .A2(new_n648), .A3(new_n805), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n814), .B2(new_n815), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n819), .A2(new_n866), .A3(new_n647), .A4(new_n813), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n864), .B1(new_n868), .B2(new_n720), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n826), .B1(new_n869), .B2(new_n598), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n870), .B2(new_n626), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n355), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n662), .A2(new_n393), .A3(new_n415), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n862), .A2(new_n872), .A3(new_n720), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n859), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n874), .B2(G141gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  AOI221_X4 g678(.A(new_n859), .B1(new_n876), .B2(new_n879), .C1(G141gat), .C2(new_n874), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  AND3_X1   g680(.A1(new_n862), .A2(new_n873), .A3(new_n872), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n689), .A2(KEYINPUT59), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT59), .B1(new_n858), .B2(new_n689), .ZN(new_n884));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n882), .A2(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n814), .A2(new_n815), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n598), .A2(new_n719), .A3(new_n805), .A4(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n869), .B2(new_n598), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n863), .B1(new_n889), .B2(new_n626), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT120), .B(new_n861), .C1(new_n890), .C2(new_n355), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n865), .B(new_n867), .C1(new_n545), .C2(new_n546), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n598), .B1(new_n893), .B2(new_n806), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n719), .A2(new_n805), .ZN(new_n895));
  INV_X1    g694(.A(new_n887), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n674), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n626), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n355), .B1(new_n898), .B2(new_n829), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n892), .B1(new_n899), .B2(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n685), .B1(new_n824), .B2(new_n826), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n453), .C1(new_n901), .C2(new_n863), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n891), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(new_n648), .A3(new_n873), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n886), .B1(new_n904), .B2(new_n905), .ZN(G1345gat));
  INV_X1    g705(.A(new_n858), .ZN(new_n907));
  INV_X1    g706(.A(G155gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n685), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n882), .A2(new_n685), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n908), .ZN(G1346gat));
  INV_X1    g710(.A(new_n304), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(new_n912), .A3(new_n598), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n882), .A2(new_n598), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n693), .A2(new_n416), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n860), .A2(new_n454), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(G169gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n720), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n727), .A2(new_n415), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n665), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n830), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n547), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT121), .Z(G1348gat));
  INV_X1    g724(.A(G176gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n922), .A2(new_n926), .A3(new_n682), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n917), .A2(new_n648), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT122), .A3(new_n926), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT122), .B1(new_n929), .B2(new_n926), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n223), .A3(new_n685), .ZN(new_n933));
  OAI21_X1  g732(.A(G183gat), .B1(new_n922), .B2(new_n626), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n225), .A3(new_n598), .ZN(new_n937));
  OAI21_X1  g736(.A(G190gat), .B1(new_n922), .B2(new_n674), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(KEYINPUT61), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(KEYINPUT61), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n920), .A2(new_n662), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n903), .A2(new_n720), .A3(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT124), .B(G197gat), .Z(new_n944));
  NOR2_X1   g743(.A1(new_n662), .A2(new_n355), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n860), .A2(new_n945), .A3(new_n916), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n720), .A2(new_n944), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n943), .A2(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n903), .A2(new_n683), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  AOI211_X1 g749(.A(G204gat), .B(new_n689), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n860), .A2(new_n945), .A3(new_n916), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n950), .A2(new_n954), .A3(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n903), .A2(new_n685), .A3(new_n942), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G211gat), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(KEYINPUT127), .A3(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n946), .A2(G211gat), .A3(new_n626), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n965), .A2(new_n969), .ZN(G1354gat));
  NAND3_X1  g769(.A1(new_n903), .A2(new_n598), .A3(new_n942), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G218gat), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n674), .A2(G218gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n946), .B2(new_n973), .ZN(G1355gat));
endmodule


