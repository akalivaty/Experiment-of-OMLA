//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n189), .A3(G143), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G146), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n189), .A2(KEYINPUT65), .A3(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n191), .B(new_n193), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n198), .A2(new_n201), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n191), .A2(new_n193), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n195), .A2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n190), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n205), .A2(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n202), .B2(new_n217), .ZN(new_n218));
  AND4_X1   g032(.A1(new_n216), .A2(new_n217), .A3(new_n190), .A4(new_n206), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n204), .B1(new_n221), .B2(G125), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G224), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT69), .B(G119), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G116), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n226), .B2(new_n227), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n230), .B(G113), .C1(new_n234), .C2(new_n229), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(new_n233), .C1(new_n227), .C2(new_n226), .ZN(new_n238));
  INV_X1    g052(.A(G104), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n239), .B2(G107), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  INV_X1    g055(.A(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G104), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(G107), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n239), .A2(G107), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n242), .A2(G104), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n238), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n234), .A2(new_n236), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n238), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n240), .A2(new_n243), .A3(new_n245), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G101), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n246), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G122), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(new_n260), .A3(new_n262), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n267), .A3(new_n263), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n225), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n235), .A2(new_n238), .A3(new_n250), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n262), .B(KEYINPUT8), .ZN(new_n271));
  INV_X1    g085(.A(new_n238), .ZN(new_n272));
  INV_X1    g086(.A(G113), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n228), .B2(new_n229), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT5), .B(new_n233), .C1(new_n226), .C2(new_n227), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n270), .B(new_n271), .C1(new_n276), .C2(new_n250), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n278));
  INV_X1    g092(.A(new_n224), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT7), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n204), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n211), .A2(new_n212), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(G128), .A3(new_n214), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n198), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n217), .A2(new_n190), .A3(new_n206), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n202), .A2(new_n216), .A3(new_n217), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(G125), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n278), .B(new_n281), .C1(new_n282), .C2(new_n290), .ZN(new_n291));
  OAI221_X1 g105(.A(new_n204), .B1(new_n280), .B2(new_n279), .C1(new_n221), .C2(G125), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n277), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n278), .B1(new_n222), .B2(new_n281), .ZN(new_n294));
  INV_X1    g108(.A(new_n265), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n269), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n269), .A2(new_n297), .A3(new_n298), .A4(new_n300), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n188), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(G234), .A2(G237), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n305), .A2(G952), .A3(new_n223), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n305), .A2(G902), .A3(G953), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT21), .B(G898), .Z(new_n310));
  OAI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G478), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT15), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G122), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n316), .A2(new_n242), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n227), .A2(KEYINPUT14), .A3(G122), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT14), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n317), .B1(new_n320), .B2(G107), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n210), .A2(G143), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n195), .A2(KEYINPUT93), .A3(G128), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT93), .B1(new_n195), .B2(G128), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT95), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT93), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n210), .B2(G143), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n195), .A2(KEYINPUT93), .A3(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT95), .A3(new_n322), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n327), .A2(new_n332), .A3(G134), .ZN(new_n333));
  AOI21_X1  g147(.A(G134), .B1(new_n327), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n321), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT97), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G134), .ZN(new_n338));
  INV_X1    g152(.A(new_n332), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT95), .B1(new_n331), .B2(new_n322), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n332), .A3(G134), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT97), .A3(new_n321), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n331), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n322), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n346), .A2(new_n331), .ZN(new_n349));
  OAI21_X1  g163(.A(G134), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n316), .B(G107), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n341), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT96), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n334), .A2(new_n351), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT96), .A3(new_n350), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT9), .B(G234), .Z(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT74), .B(G217), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n223), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n345), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n345), .B2(new_n358), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n298), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT98), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n335), .A2(new_n336), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT97), .B1(new_n343), .B2(new_n321), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT96), .B1(new_n356), .B2(new_n350), .ZN(new_n369));
  AND4_X1   g183(.A1(KEYINPUT96), .A2(new_n350), .A3(new_n341), .A4(new_n352), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n361), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n345), .A2(new_n358), .A3(new_n362), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT98), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n298), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n315), .B1(new_n366), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n314), .B1(new_n365), .B2(KEYINPUT98), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT99), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n375), .B1(new_n374), .B2(new_n298), .ZN(new_n380));
  AOI211_X1 g194(.A(KEYINPUT98), .B(G902), .C1(new_n372), .C2(new_n373), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n314), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT99), .ZN(new_n383));
  INV_X1    g197(.A(new_n378), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n312), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G469), .ZN(new_n387));
  XOR2_X1   g201(.A(G110), .B(G140), .Z(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT81), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n223), .A2(G227), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n210), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(new_n202), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n250), .B1(new_n289), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI211_X1 g211(.A(KEYINPUT82), .B(new_n250), .C1(new_n289), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n203), .A2(new_n257), .A3(new_n259), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n285), .A2(new_n289), .A3(KEYINPUT70), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT70), .B1(new_n285), .B2(new_n289), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT10), .B(new_n251), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT85), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT11), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n406), .A2(new_n407), .B1(new_n338), .B2(G137), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n406), .A2(new_n407), .B1(new_n338), .B2(G137), .ZN(new_n409));
  INV_X1    g223(.A(G137), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G131), .ZN(new_n413));
  INV_X1    g227(.A(G131), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n408), .A2(new_n409), .A3(new_n414), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n399), .A2(new_n417), .A3(new_n400), .A4(new_n403), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n405), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n416), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n399), .A2(new_n420), .A3(new_n400), .A4(new_n403), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n391), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n221), .A2(new_n250), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n397), .B2(new_n398), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n426), .B2(new_n416), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n426), .A2(KEYINPUT83), .A3(new_n423), .A4(new_n416), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n391), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n387), .B(new_n298), .C1(new_n422), .C2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n387), .A2(new_n298), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n391), .ZN(new_n437));
  INV_X1    g251(.A(new_n421), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n431), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n421), .A2(new_n441), .A3(new_n391), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n419), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n443), .A3(G469), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n434), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G221), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n359), .B2(new_n298), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OR2_X1    g264(.A1(KEYINPUT71), .A2(G237), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT71), .A2(G237), .ZN(new_n452));
  AOI21_X1  g266(.A(G953), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(G143), .B1(new_n453), .B2(G214), .ZN(new_n454));
  AND2_X1   g268(.A1(KEYINPUT71), .A2(G237), .ZN(new_n455));
  NOR2_X1   g269(.A1(KEYINPUT71), .A2(G237), .ZN(new_n456));
  OAI211_X1 g270(.A(G214), .B(new_n223), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n195), .ZN(new_n458));
  OAI21_X1  g272(.A(G131), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n195), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n451), .A2(new_n452), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(G143), .A3(G214), .A4(new_n223), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n463), .A3(new_n414), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT16), .ZN(new_n466));
  INV_X1    g280(.A(G140), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(G125), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT77), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(G125), .ZN(new_n470));
  INV_X1    g284(.A(G125), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G140), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(KEYINPUT76), .A3(new_n466), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n475));
  XNOR2_X1  g289(.A(G125), .B(G140), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(KEYINPUT16), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n469), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n189), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n469), .B(G146), .C1(new_n474), .C2(new_n477), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n414), .B1(new_n461), .B2(new_n463), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT17), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n465), .A2(new_n479), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n461), .B(new_n463), .C1(new_n484), .C2(new_n414), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n476), .A2(KEYINPUT79), .A3(new_n189), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT79), .B1(new_n476), .B2(new_n189), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n486), .A2(new_n487), .B1(new_n189), .B2(new_n476), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n485), .B(new_n488), .C1(new_n459), .C2(new_n484), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT88), .B(G104), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT89), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n483), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n476), .B(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n189), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n461), .A2(new_n463), .A3(new_n414), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n480), .B(new_n496), .C1(new_n497), .C2(new_n481), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n492), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  NOR2_X1   g317(.A1(G475), .A2(G902), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n502), .B2(new_n504), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n502), .A2(KEYINPUT90), .A3(new_n503), .A4(new_n504), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT91), .B(G475), .Z(new_n511));
  AND2_X1   g325(.A1(new_n483), .A2(new_n489), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n494), .B1(new_n512), .B2(new_n492), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n513), .B2(new_n298), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(KEYINPUT92), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n386), .A2(new_n450), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n416), .A2(new_n203), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n215), .B2(new_n220), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n285), .A2(new_n289), .A3(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n410), .A2(G134), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n338), .A2(G137), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n415), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n524), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n254), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT28), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n537), .A3(new_n534), .ZN(new_n538));
  INV_X1    g352(.A(new_n533), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n536), .A2(new_n538), .B1(new_n254), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n453), .A2(G210), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(G101), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n532), .B1(new_n401), .B2(new_n402), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n523), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n532), .B1(new_n215), .B2(new_n220), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n523), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT30), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n254), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n555), .A2(new_n535), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n544), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n254), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n537), .B1(new_n533), .B2(new_n534), .ZN(new_n559));
  AND4_X1   g373(.A1(new_n537), .A2(new_n550), .A3(new_n534), .A4(new_n523), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n546), .B1(new_n561), .B2(new_n545), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n548), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n555), .A2(new_n535), .A3(new_n544), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT31), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n545), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n568));
  NAND4_X1  g382(.A1(new_n555), .A2(new_n535), .A3(new_n544), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G472), .A2(G902), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT32), .B1(new_n572), .B2(KEYINPUT73), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n574), .B(new_n575), .C1(new_n570), .C2(new_n571), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n564), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  INV_X1    g392(.A(G234), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n446), .A2(new_n579), .A3(G953), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n578), .B(new_n580), .Z(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT23), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT69), .B(G119), .Z(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(G128), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G110), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n210), .A2(G119), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(KEYINPUT75), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT24), .B(G110), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n593), .B(new_n594), .C1(KEYINPUT75), .C2(new_n586), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n486), .A2(new_n487), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n480), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n591), .B1(new_n590), .B2(new_n595), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n588), .A2(new_n589), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n479), .A2(new_n480), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n593), .B1(KEYINPUT75), .B2(new_n586), .ZN(new_n603));
  INV_X1    g417(.A(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n582), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  OR2_X1    g422(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n606), .B(new_n581), .C1(new_n598), .C2(new_n599), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n608), .A2(new_n298), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n360), .B1(new_n579), .B2(G902), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n608), .ZN(new_n616));
  INV_X1    g430(.A(new_n610), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n615), .A2(G902), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n613), .A2(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n577), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n522), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  INV_X1    g437(.A(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n570), .A2(new_n298), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n572), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n624), .A2(new_n449), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n311), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n188), .B(new_n629), .C1(new_n302), .C2(new_n303), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n363), .B2(new_n364), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n372), .A2(KEYINPUT33), .A3(new_n373), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n313), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n365), .A2(G478), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n313), .A2(new_n298), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT92), .B1(new_n510), .B2(new_n515), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n517), .B(new_n514), .C1(new_n508), .C2(new_n509), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n630), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n628), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AND2_X1   g458(.A1(new_n379), .A2(new_n385), .ZN(new_n645));
  INV_X1    g459(.A(new_n506), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n514), .B1(new_n505), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n645), .A2(new_n630), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n628), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND2_X1  g465(.A1(new_n613), .A2(new_n615), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n600), .A2(new_n607), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n582), .A2(KEYINPUT36), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n619), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n522), .A2(new_n572), .A3(new_n626), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G12));
  OAI21_X1  g475(.A(new_n307), .B1(new_n309), .B2(G900), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n379), .A2(new_n385), .A3(new_n647), .A4(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n445), .A2(new_n448), .A3(new_n304), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n577), .A3(new_n664), .A4(new_n657), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XOR2_X1   g480(.A(new_n662), .B(KEYINPUT39), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n450), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n188), .A4(new_n657), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n556), .A2(new_n545), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n535), .A2(new_n545), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n533), .A2(new_n534), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n298), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n573), .B2(new_n576), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n680), .B(new_n677), .C1(new_n573), .C2(new_n576), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n379), .B(new_n385), .C1(new_n638), .C2(new_n639), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n302), .A2(new_n303), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n672), .A2(new_n682), .A3(new_n684), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  OAI211_X1 g503(.A(new_n637), .B(new_n662), .C1(new_n638), .C2(new_n639), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n577), .A3(new_n664), .A4(new_n657), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  OAI21_X1  g507(.A(new_n298), .B1(new_n422), .B2(new_n433), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n448), .A3(new_n434), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n641), .A2(new_n577), .A3(new_n620), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND3_X1  g514(.A1(new_n648), .A2(new_n621), .A3(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NAND4_X1  g516(.A1(new_n577), .A2(new_n386), .A3(new_n521), .A4(new_n657), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n696), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n231), .ZN(G21));
  INV_X1    g519(.A(new_n304), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT104), .B1(new_n683), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n645), .A2(new_n708), .A3(new_n520), .A4(new_n304), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n566), .B(new_n569), .C1(new_n544), .C2(new_n540), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(new_n571), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n626), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n625), .A2(KEYINPUT103), .A3(G472), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n620), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n696), .A2(new_n629), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n710), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NOR2_X1   g535(.A1(new_n690), .A2(new_n696), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n716), .A3(new_n304), .A4(new_n657), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT105), .B(G125), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G27));
  NOR2_X1   g539(.A1(new_n685), .A2(new_n188), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n449), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n691), .A3(new_n577), .A4(new_n620), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n570), .A2(new_n575), .A3(new_n571), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n575), .B1(new_n570), .B2(new_n571), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n564), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n620), .A3(KEYINPUT42), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n520), .A2(new_n637), .A3(new_n662), .A4(new_n726), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT106), .B1(new_n737), .B2(new_n450), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n735), .A2(new_n736), .A3(new_n739), .A4(new_n449), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n731), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(new_n731), .C1(new_n738), .C2(new_n740), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND2_X1  g560(.A1(new_n621), .A2(new_n728), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n663), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(new_n637), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n520), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n627), .A3(new_n657), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n727), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n439), .A2(new_n443), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n435), .B1(new_n758), .B2(G469), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n434), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n762), .A2(new_n448), .A3(new_n668), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n756), .B(new_n763), .C1(new_n755), .C2(new_n754), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n762), .B2(new_n448), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n762), .A2(new_n766), .A3(new_n448), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n577), .A2(new_n620), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n770), .A2(new_n736), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  AND3_X1   g587(.A1(new_n753), .A2(new_n306), .A3(new_n718), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n697), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n687), .A2(new_n187), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n716), .A2(new_n657), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n697), .A2(new_n726), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT117), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(KEYINPUT117), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n307), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n753), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n777), .A2(KEYINPUT50), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n682), .A2(new_n624), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n521), .A3(new_n751), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n785), .B(new_n788), .C1(KEYINPUT50), .C2(new_n777), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(KEYINPUT118), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n695), .A2(new_n447), .A3(new_n434), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT116), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n774), .A2(new_n726), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(KEYINPUT51), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n798), .B1(new_n770), .B2(new_n795), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n789), .B2(new_n801), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n792), .A2(new_n799), .B1(new_n802), .B2(new_n790), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  INV_X1    g618(.A(new_n749), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n742), .B2(new_n744), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n698), .B1(new_n703), .B2(new_n696), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n720), .A3(new_n701), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT108), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n808), .A2(new_n720), .A3(new_n811), .A4(new_n701), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n716), .A2(new_n520), .A3(new_n637), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n377), .A2(new_n378), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n577), .A2(new_n815), .A3(new_n647), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n657), .A3(new_n662), .A4(new_n728), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n520), .A2(new_n637), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT109), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n819), .B(KEYINPUT109), .C1(new_n520), .C2(new_n815), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n628), .A4(new_n630), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n818), .A2(new_n622), .A3(new_n658), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n806), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n657), .B1(new_n679), .B2(new_n681), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n710), .A3(new_n450), .A4(new_n662), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n723), .A2(new_n665), .A3(new_n692), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n828), .A2(KEYINPUT52), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n826), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n829), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(KEYINPUT113), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n825), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(KEYINPUT110), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n828), .A2(new_n829), .A3(new_n841), .A4(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n723), .A2(new_n665), .A3(new_n692), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n449), .B1(new_n707), .B2(new_n709), .ZN(new_n847));
  INV_X1    g661(.A(new_n662), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n657), .B(new_n848), .C1(new_n679), .C2(new_n681), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n845), .B1(new_n850), .B2(KEYINPUT52), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n833), .A2(KEYINPUT111), .A3(new_n834), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n843), .A2(new_n844), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n831), .A2(KEYINPUT111), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n845), .B(KEYINPUT52), .C1(new_n828), .C2(new_n829), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n844), .B1(new_n857), .B2(new_n843), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n806), .A2(new_n813), .A3(new_n824), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n804), .ZN(new_n861));
  OAI221_X1 g675(.A(KEYINPUT54), .B1(new_n804), .B2(new_n839), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n809), .A2(KEYINPUT114), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n823), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n804), .B1(new_n809), .B2(KEYINPUT114), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n741), .A3(new_n749), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n841), .B1(new_n850), .B2(KEYINPUT52), .ZN(new_n867));
  INV_X1    g681(.A(new_n842), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n851), .A2(new_n852), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT112), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n866), .B1(new_n871), .B2(new_n853), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n832), .A2(new_n837), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n860), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n787), .ZN(new_n877));
  OAI211_X1 g691(.A(G952), .B(new_n223), .C1(new_n877), .C2(new_n819), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n304), .B2(new_n775), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n803), .A2(new_n862), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n734), .A2(new_n620), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n784), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  OAI22_X1  g697(.A1(new_n880), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n695), .A2(new_n434), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(KEYINPUT49), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n448), .B1(new_n885), .B2(KEYINPUT49), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n188), .A4(new_n687), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n786), .A2(new_n752), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n223), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n866), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n854), .B2(new_n858), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n804), .B1(new_n825), .B2(new_n838), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n298), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G210), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n266), .A2(new_n268), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n225), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  INV_X1    g719(.A(new_n904), .ZN(new_n906));
  AOI211_X1 g720(.A(KEYINPUT119), .B(new_n906), .C1(new_n897), .C2(new_n898), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(G51));
  XOR2_X1   g722(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n435), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n909), .A2(new_n435), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n894), .B2(new_n895), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n910), .B(new_n911), .C1(new_n913), .C2(new_n875), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n422), .B2(new_n433), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n896), .A2(G469), .A3(new_n758), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n891), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n892), .B1(new_n919), .B2(new_n502), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT121), .B1(new_n919), .B2(new_n502), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  INV_X1    g736(.A(new_n502), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(G60));
  AND2_X1   g739(.A1(new_n632), .A2(new_n633), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n636), .B(KEYINPUT59), .Z(new_n927));
  OAI211_X1 g741(.A(new_n926), .B(new_n927), .C1(new_n913), .C2(new_n875), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n928), .A2(KEYINPUT122), .A3(new_n892), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT122), .B1(new_n928), .B2(new_n892), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n876), .A2(new_n862), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n926), .B1(new_n931), .B2(new_n927), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n894), .B2(new_n895), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n655), .ZN(new_n937));
  INV_X1    g751(.A(new_n935), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n872), .B2(new_n874), .ZN(new_n939));
  INV_X1    g753(.A(new_n618), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n892), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n939), .A2(new_n945), .A3(new_n940), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n939), .B2(new_n940), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n892), .A2(KEYINPUT61), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n936), .B2(new_n655), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT124), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n941), .A2(KEYINPUT123), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n939), .A2(new_n945), .A3(new_n940), .ZN(new_n953));
  AND4_X1   g767(.A1(KEYINPUT124), .A2(new_n952), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n944), .B1(new_n951), .B2(new_n954), .ZN(G66));
  AOI21_X1  g769(.A(new_n223), .B1(new_n310), .B2(G224), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n813), .A2(new_n622), .A3(new_n658), .A4(new_n822), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n223), .ZN(new_n958));
  INV_X1    g772(.A(G898), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n902), .B1(new_n959), .B2(G953), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  NAND2_X1  g775(.A1(new_n688), .A2(new_n829), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NAND4_X1  g777(.A1(new_n748), .A2(new_n668), .A3(new_n821), .A4(new_n820), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n764), .A3(new_n772), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n223), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n551), .A2(new_n554), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(new_n495), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  NAND2_X1  g784(.A1(G900), .A2(G953), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n763), .A2(new_n710), .A3(new_n881), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n806), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n764), .A3(new_n772), .A4(new_n829), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n970), .B(new_n971), .C1(new_n974), .C2(G953), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n966), .A2(KEYINPUT125), .A3(new_n968), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT125), .B1(new_n966), .B2(new_n968), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n977), .B(KEYINPUT126), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n965), .B2(new_n957), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n673), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n974), .B2(new_n957), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n545), .A3(new_n556), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n892), .A3(new_n989), .ZN(new_n990));
  OAI22_X1  g804(.A1(new_n859), .A2(new_n861), .B1(new_n804), .B2(new_n839), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT127), .B1(new_n556), .B2(new_n544), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(new_n557), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n985), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n992), .B2(new_n995), .ZN(G57));
endmodule


