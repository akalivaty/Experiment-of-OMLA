//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n452, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G234));
  INV_X1    g026(.A(G2106), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  OAI22_X1  g035(.A1(new_n456), .A2(new_n452), .B1(new_n449), .B2(new_n457), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g056(.A1(new_n471), .A2(new_n478), .A3(new_n481), .ZN(G160));
  NAND4_X1  g057(.A1(new_n476), .A2(new_n472), .A3(new_n474), .A4(new_n466), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n474), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n476), .A2(new_n472), .A3(G2105), .A4(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT71), .A3(G124), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  INV_X1    g066(.A(G124), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n490), .B2(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n476), .A2(new_n472), .A3(new_n496), .A4(new_n466), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(G138), .A3(new_n474), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n464), .A2(new_n466), .ZN(new_n502));
  AOI22_X1  g077(.A1(KEYINPUT4), .A2(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n474), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n488), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(new_n513), .A3(G62), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n510), .B1(new_n517), .B2(new_n516), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n515), .A2(new_n524), .ZN(G166));
  NAND2_X1  g100(.A1(new_n520), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT5), .B(G543), .Z(new_n530));
  OR2_X1    g105(.A1(new_n516), .A2(new_n517), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n509), .B1(new_n538), .B2(KEYINPUT74), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(KEYINPUT74), .B2(new_n538), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n530), .A2(new_n518), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n541), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n520), .A2(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n544), .B(new_n545), .C1(new_n509), .C2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT75), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n523), .A2(KEYINPUT77), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT77), .B1(new_n523), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(KEYINPUT76), .A2(G53), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n531), .A2(G543), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n520), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n530), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n561), .A2(new_n563), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n558), .A2(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(G171), .A2(KEYINPUT78), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n540), .A2(new_n542), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND2_X1  g151(.A1(new_n541), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n520), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n509), .ZN(new_n582));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n523), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  INV_X1    g163(.A(G72), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n530), .A2(new_n588), .B1(new_n589), .B2(new_n519), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT79), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n592), .B1(new_n589), .B2(new_n519), .C1(new_n530), .C2(new_n588), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(G651), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n541), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G290));
  AND3_X1   g174(.A1(new_n531), .A2(G92), .A3(new_n510), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n530), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n573), .B2(G868), .ZN(G284));
  XNOR2_X1  g183(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  AND2_X1   g188(.A1(new_n601), .A2(new_n605), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(new_n483), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G135), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT82), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n489), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n474), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT83), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n502), .A2(new_n479), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(KEYINPUT13), .B(G2100), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n644), .A2(new_n647), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  INV_X1    g249(.A(new_n669), .ZN(new_n675));
  INV_X1    g250(.A(new_n672), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n674), .B(new_n678), .C1(new_n675), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  NOR2_X1   g260(.A1(G6), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n586), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT32), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1981), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G22), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G166), .B2(G16), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n691), .A2(G1971), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(G1971), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  NOR4_X1   g274(.A1(new_n689), .A2(new_n692), .A3(new_n693), .A4(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n694), .A2(G24), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G290), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  INV_X1    g284(.A(G119), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n488), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT88), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(G107), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G2105), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n621), .A2(G131), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(new_n708), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n702), .A2(new_n703), .A3(new_n707), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT36), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n549), .A2(new_n694), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n694), .B2(G19), .ZN(new_n724));
  INV_X1    g299(.A(G1341), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G160), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2084), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n724), .A2(new_n725), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n694), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n694), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1961), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n726), .A2(new_n733), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n708), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G105), .B2(new_n479), .ZN(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n488), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n621), .B2(G141), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n708), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT93), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n738), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n708), .A2(G26), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n757));
  INV_X1    g332(.A(G140), .ZN(new_n758));
  INV_X1    g333(.A(G128), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n757), .B1(new_n483), .B2(new_n758), .C1(new_n759), .C2(new_n488), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n762), .A2(KEYINPUT91), .A3(G29), .ZN(new_n763));
  AOI21_X1  g338(.A(KEYINPUT91), .B1(new_n762), .B2(G29), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G4), .A2(G16), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n614), .B2(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G1348), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n474), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G139), .B2(new_n621), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(new_n708), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n708), .B2(G33), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n770), .B1(new_n779), .B2(G2072), .ZN(new_n780));
  INV_X1    g355(.A(G2072), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n778), .A2(new_n781), .B1(G1348), .B2(new_n769), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT99), .B(KEYINPUT23), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n694), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n708), .A2(G27), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G164), .B2(new_n708), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT97), .B(G2078), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n780), .A2(new_n782), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n753), .A2(new_n767), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n736), .A2(G1961), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT95), .Z(new_n796));
  OR2_X1    g371(.A1(new_n628), .A2(new_n708), .ZN(new_n797));
  NOR2_X1   g372(.A1(G168), .A2(new_n694), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n694), .B2(G21), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(G28), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n708), .B1(new_n803), .B2(G28), .ZN(new_n805));
  AND2_X1   g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  NOR2_X1   g381(.A1(KEYINPUT31), .A2(G11), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n799), .B2(new_n800), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n796), .A2(new_n797), .A3(new_n802), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G35), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G162), .B2(G29), .ZN(new_n813));
  INV_X1    g388(.A(G2090), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n794), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n722), .A2(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  AOI22_X1  g395(.A1(new_n541), .A2(G93), .B1(new_n520), .B2(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n509), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NOR2_X1   g400(.A1(new_n606), .A2(new_n615), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n823), .A2(new_n547), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n548), .B2(new_n823), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n828), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT101), .Z(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n832), .B2(new_n833), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n825), .B1(new_n835), .B2(new_n837), .ZN(G145));
  INV_X1    g413(.A(G37), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n717), .B(new_n631), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n621), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n489), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n474), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n840), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n762), .B(G164), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n747), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n776), .B(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n776), .A2(new_n852), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n846), .B1(new_n854), .B2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n628), .B(new_n731), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n847), .B(new_n848), .C1(new_n854), .C2(new_n856), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n839), .B(new_n862), .C1(new_n864), .C2(new_n861), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g441(.A(G290), .B(G305), .ZN(new_n867));
  XNOR2_X1  g442(.A(G166), .B(G288), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT42), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n617), .B(KEYINPUT104), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n831), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n614), .B2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n614), .A2(G299), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n611), .A2(new_n606), .A3(KEYINPUT105), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n880), .B1(new_n874), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n872), .B(new_n888), .ZN(new_n889));
  MUX2_X1   g464(.A(new_n823), .B(new_n889), .S(G868), .Z(G295));
  MUX2_X1   g465(.A(new_n823), .B(new_n889), .S(G868), .Z(G331));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  INV_X1    g467(.A(new_n869), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n573), .A2(G168), .ZN(new_n894));
  NOR2_X1   g469(.A1(G171), .A2(G168), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n830), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G286), .B1(new_n569), .B2(new_n572), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n831), .B1(new_n898), .B2(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n899), .A3(KEYINPUT108), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n894), .A2(new_n901), .A3(new_n830), .A4(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n882), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n879), .A2(KEYINPUT41), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(KEYINPUT109), .A3(new_n884), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n897), .A2(new_n899), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n906), .B(new_n907), .C1(KEYINPUT109), .C2(new_n905), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n893), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n897), .A2(new_n899), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n882), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n881), .A2(new_n884), .A3(new_n886), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n893), .B(new_n912), .C1(new_n903), .C2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n910), .A2(new_n914), .A3(new_n915), .A4(new_n839), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n839), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT110), .B1(new_n917), .B2(new_n909), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n892), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n912), .B1(new_n903), .B2(new_n913), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n869), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT44), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n910), .A2(new_n892), .A3(new_n839), .A4(new_n914), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n921), .B2(new_n892), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(KEYINPUT127), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT125), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT116), .ZN(new_n931));
  INV_X1    g506(.A(G1981), .ZN(new_n932));
  INV_X1    g507(.A(new_n582), .ZN(new_n933));
  INV_X1    g508(.A(new_n585), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n582), .A2(new_n585), .A3(G1981), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT49), .ZN(new_n938));
  INV_X1    g513(.A(G8), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n505), .A2(new_n506), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n489), .B2(G126), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n501), .A2(new_n502), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G1384), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AND4_X1   g520(.A1(G40), .A2(new_n470), .A3(new_n477), .A4(new_n480), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n939), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT49), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n931), .B(new_n948), .C1(new_n935), .C2(new_n936), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1976), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n951), .B2(G288), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT52), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(G288), .B2(new_n951), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n947), .B(new_n954), .C1(new_n951), .C2(G288), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(G1971), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n503), .B2(new_n507), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT45), .B(new_n958), .C1(new_n503), .C2(new_n507), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n946), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n959), .B2(new_n961), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(new_n958), .C1(new_n503), .C2(new_n507), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n967), .A2(new_n969), .A3(new_n946), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n814), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(G166), .B2(new_n939), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT55), .B(G8), .C1(new_n515), .C2(new_n524), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n956), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(KEYINPUT114), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n966), .A2(new_n971), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n975), .A2(new_n982), .A3(new_n976), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n975), .B2(new_n976), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n979), .A2(G8), .A3(new_n981), .A4(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT123), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n978), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n978), .B2(new_n986), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n959), .A2(new_n961), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n470), .A2(new_n477), .A3(G40), .A4(new_n480), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n945), .B2(KEYINPUT45), .ZN(new_n994));
  INV_X1    g569(.A(G2078), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n962), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n945), .A2(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n963), .A2(new_n946), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n997), .A2(G2078), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n967), .A2(new_n969), .A3(new_n946), .ZN(new_n1003));
  INV_X1    g578(.A(G1961), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1001), .A2(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n573), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n800), .B1(new_n999), .B2(new_n1000), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n993), .B1(new_n959), .B2(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(G2084), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n969), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(G168), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G286), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(G8), .A3(new_n1012), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1017), .B2(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1007), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n930), .B1(new_n990), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n978), .A2(new_n986), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT123), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n978), .A2(new_n986), .A3(new_n987), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1020), .A3(new_n930), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1014), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT126), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(KEYINPUT62), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT126), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n929), .B1(new_n1021), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n992), .A2(new_n994), .A3(new_n962), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1035), .A2(new_n957), .B1(new_n970), .B2(new_n814), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n1036), .B2(new_n980), .ZN(new_n1037));
  INV_X1    g612(.A(new_n981), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n977), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n939), .B(G286), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT63), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n956), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1039), .A2(new_n986), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n978), .A2(new_n986), .A3(new_n1040), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT63), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n986), .A2(new_n956), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n950), .A2(new_n951), .A3(new_n696), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(G1981), .B2(G305), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n947), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n558), .A2(new_n567), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n558), .B2(new_n567), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n992), .A2(new_n994), .A3(new_n962), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1003), .A2(new_n787), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n959), .A2(new_n993), .A3(G2067), .ZN(new_n1059));
  INV_X1    g634(.A(G1348), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1003), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1058), .B1(new_n1061), .B2(new_n606), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1348), .B1(new_n1009), .B2(new_n969), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT118), .B(new_n614), .C1(new_n1063), .C2(new_n1059), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1055), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1057), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR4_X1   g642(.A1(new_n1063), .A2(KEYINPUT60), .A3(new_n606), .A4(new_n1059), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1061), .B2(new_n614), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n606), .B1(new_n1063), .B2(new_n1059), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n945), .A2(new_n946), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT119), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT119), .B(new_n1075), .C1(new_n959), .C2(new_n993), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1996), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n992), .A2(new_n994), .A3(new_n1080), .A4(new_n962), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1073), .B1(new_n1082), .B2(new_n549), .ZN(new_n1083));
  AOI211_X1 g658(.A(KEYINPUT59), .B(new_n548), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1072), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1055), .A2(new_n1053), .A3(new_n1056), .A4(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1067), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n991), .A2(new_n963), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1002), .B1(new_n946), .B2(KEYINPUT122), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n993), .A2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n997), .B2(new_n996), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT121), .B1(new_n970), .B2(G1961), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1003), .A2(new_n1098), .A3(new_n1004), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1100), .A3(G301), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1007), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n998), .A2(new_n1005), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1105), .B2(G301), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1106), .A2(new_n1108), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1090), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1045), .B(new_n1049), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1023), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT125), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1116), .A2(KEYINPUT127), .A3(new_n1025), .A4(new_n1032), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1104), .A2(new_n1118), .A3(new_n1028), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n990), .A2(new_n1119), .A3(new_n1090), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(KEYINPUT124), .A3(new_n1045), .A4(new_n1049), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1034), .A2(new_n1114), .A3(new_n1117), .A4(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n991), .A2(new_n993), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(G1996), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n747), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT111), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n762), .B(new_n766), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1080), .B2(new_n747), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n717), .A2(new_n719), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n717), .A2(new_n719), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1123), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(G290), .B(G1986), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n1123), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1122), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1125), .B(KEYINPUT46), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1124), .B1(new_n1128), .B2(new_n747), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT47), .Z(new_n1141));
  NOR3_X1   g716(.A1(G290), .A2(new_n1124), .A3(G1986), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT48), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1134), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n762), .A2(G2067), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1124), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1137), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g724(.A(G319), .B1(new_n649), .B2(new_n650), .ZN(new_n1151));
  NOR3_X1   g725(.A1(G229), .A2(G227), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n865), .A3(new_n1152), .ZN(G225));
  INV_X1    g727(.A(G225), .ZN(G308));
endmodule


