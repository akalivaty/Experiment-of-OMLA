//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G137), .ZN(new_n461));
  INV_X1    g036(.A(G101), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G2104), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n458), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT66), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  AND2_X1   g045(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n459), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n459), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n460), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n459), .A2(KEYINPUT4), .A3(G138), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(new_n459), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n459), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n488), .A2(new_n458), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n497), .B2(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n495), .A3(KEYINPUT6), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(G88), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n498), .A2(new_n500), .ZN(new_n508));
  INV_X1    g083(.A(new_n496), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G543), .A3(new_n509), .ZN(new_n510));
  OAI221_X1 g085(.A(new_n505), .B1(new_n506), .B2(new_n495), .C1(new_n507), .C2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  AOI211_X1 g088(.A(new_n513), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n504), .A2(KEYINPUT69), .A3(G63), .A4(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n514), .A2(G51), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT70), .A2(G89), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT70), .A2(G89), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n508), .A2(new_n509), .A3(new_n504), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n527), .B1(new_n526), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n522), .B1(new_n530), .B2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n502), .B2(new_n503), .ZN(new_n535));
  AND2_X1   g110(.A1(G77), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n508), .A2(G90), .A3(new_n509), .A4(new_n504), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n508), .A2(G52), .A3(G543), .A4(new_n509), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G171));
  NAND3_X1  g115(.A1(new_n501), .A2(G81), .A3(new_n504), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n501), .A2(G43), .A3(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n502), .B2(new_n503), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  AND3_X1   g128(.A1(new_n501), .A2(G91), .A3(new_n504), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n504), .B2(G65), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n495), .B1(new_n557), .B2(KEYINPUT74), .ZN(new_n558));
  OAI21_X1  g133(.A(G65), .B1(new_n517), .B2(new_n518), .ZN(new_n559));
  AOI21_X1  g134(.A(KEYINPUT74), .B1(new_n559), .B2(new_n555), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n554), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G53), .A2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n501), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT73), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n509), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n501), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n562), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND4_X1  g150(.A1(new_n508), .A2(G87), .A3(new_n509), .A4(new_n504), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n510), .C2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n514), .A2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n501), .A2(G86), .A3(new_n504), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n519), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(G305));
  NAND3_X1  g161(.A1(new_n501), .A2(G85), .A3(new_n504), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n501), .A2(G47), .A3(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n502), .B2(new_n503), .ZN(new_n590));
  AND2_X1   g165(.A1(G72), .A2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n502), .B2(new_n503), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(KEYINPUT75), .A2(G79), .A3(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n508), .A2(G54), .A3(G543), .A4(new_n509), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n508), .A2(G92), .A3(new_n509), .A4(new_n504), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n501), .A2(KEYINPUT10), .A3(G92), .A4(new_n504), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n594), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n594), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n501), .A2(G91), .A3(new_n504), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n559), .A2(KEYINPUT74), .A3(new_n555), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n560), .ZN(new_n616));
  INV_X1    g191(.A(new_n572), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n571), .B1(new_n501), .B2(new_n566), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n619), .B2(new_n570), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n612), .B1(G868), .B2(new_n620), .ZN(G297));
  OAI21_X1  g196(.A(new_n612), .B1(G868), .B2(new_n620), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n609), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g203(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n631), .A2(new_n632), .B1(KEYINPUT76), .B2(G2100), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  OR3_X1    g209(.A1(new_n634), .A2(KEYINPUT76), .A3(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n474), .A2(G123), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n477), .A2(G135), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n634), .B1(KEYINPUT76), .B2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(G2096), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n635), .A2(new_n641), .A3(new_n642), .A4(new_n643), .ZN(G156));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT77), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n653), .B2(new_n654), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT78), .Z(new_n663));
  AOI21_X1  g238(.A(new_n645), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n665), .A3(new_n660), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g247(.A(KEYINPUT80), .B(new_n664), .C1(new_n668), .C2(new_n669), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT81), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n678), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2084), .B(G2090), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n677), .B(KEYINPUT17), .Z(new_n682));
  INV_X1    g257(.A(new_n675), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n681), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n677), .A2(new_n675), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT18), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2096), .B(G2100), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n701), .B(new_n700), .S(new_n693), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1991), .B(G1996), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n704), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n703), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n706), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n707), .B2(new_n711), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1971), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n716), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G6), .A2(G16), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n719), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT85), .B(KEYINPUT34), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(G25), .A2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n474), .A2(G119), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n477), .A2(G131), .ZN(new_n736));
  OR2_X1    g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT84), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(KEYINPUT84), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n734), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  AND2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G290), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G16), .B2(G24), .ZN(new_n753));
  INV_X1    g328(.A(G1986), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(KEYINPUT87), .A3(new_n756), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n733), .A2(new_n749), .A3(new_n750), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n730), .A2(new_n732), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT86), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n760), .A3(KEYINPUT36), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n469), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT92), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G2084), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n716), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n609), .B2(new_n716), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n768), .A2(G2084), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n716), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n716), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G1961), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n548), .A2(new_n716), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n716), .B2(G19), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT88), .B(G1341), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n774), .A2(new_n775), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G168), .A2(G16), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n785), .B(new_n786), .C1(G16), .C2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT96), .B(G1966), .Z(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n746), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT28), .ZN(new_n794));
  NOR2_X1   g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT89), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n474), .B2(G128), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n477), .A2(G140), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G29), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(KEYINPUT90), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(KEYINPUT90), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n794), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2067), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n746), .A2(G33), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n458), .A2(G127), .ZN(new_n809));
  AND2_X1   g384(.A1(G115), .A2(G2104), .ZN(new_n810));
  OAI21_X1  g385(.A(G2105), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n477), .A2(G139), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT25), .Z(new_n815));
  AND3_X1   g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n808), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G2072), .Z(new_n820));
  AND2_X1   g395(.A1(new_n788), .A2(new_n790), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n807), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n477), .A2(KEYINPUT93), .A3(G141), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n824));
  INV_X1    g399(.A(G141), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n476), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT26), .Z(new_n829));
  INV_X1    g404(.A(G105), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n463), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n474), .B2(G129), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n833), .A2(KEYINPUT94), .A3(new_n746), .ZN(new_n834));
  OR2_X1    g409(.A1(G29), .A2(G32), .ZN(new_n835));
  OAI211_X1 g410(.A(KEYINPUT94), .B(new_n835), .C1(new_n833), .C2(new_n746), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT27), .B(G1996), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n746), .A2(G35), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G162), .B2(new_n746), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT29), .B(G2090), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(new_n781), .B2(new_n782), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT31), .B(G11), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT97), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT30), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(G28), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n746), .B1(new_n846), .B2(G28), .ZN(new_n848));
  OAI221_X1 g423(.A(new_n845), .B1(new_n847), .B2(new_n848), .C1(new_n640), .C2(new_n746), .ZN(new_n849));
  NOR2_X1   g424(.A1(G27), .A2(G29), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G164), .B2(G29), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G2078), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n843), .B(new_n853), .C1(new_n841), .C2(new_n842), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n716), .A2(G20), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT23), .Z(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G299), .B2(G16), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT99), .B(G1956), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT100), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n839), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n784), .A2(new_n792), .A3(new_n822), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT36), .B1(new_n758), .B2(new_n760), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n762), .A2(new_n862), .A3(new_n863), .ZN(G311));
  OR3_X1    g439(.A1(new_n762), .A2(new_n862), .A3(new_n863), .ZN(G150));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n502), .B2(new_n503), .ZN(new_n867));
  AND2_X1   g442(.A1(G80), .A2(G543), .ZN(new_n868));
  OAI21_X1  g443(.A(G651), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n508), .A2(G93), .A3(new_n509), .A4(new_n504), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n508), .A2(G55), .A3(G543), .A4(new_n509), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(KEYINPUT101), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n548), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n547), .A2(new_n872), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n607), .A2(new_n608), .ZN(new_n880));
  INV_X1    g455(.A(new_n604), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n623), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n879), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g460(.A(G860), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n874), .A2(new_n875), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G860), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT37), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(G145));
  XNOR2_X1  g466(.A(new_n469), .B(new_n640), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n481), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n802), .A2(new_n493), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n800), .A2(G164), .A3(new_n801), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n745), .B(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n818), .A2(new_n833), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n901));
  INV_X1    g476(.A(G118), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(G2105), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n477), .B2(G142), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n474), .A2(new_n905), .A3(G130), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n474), .B2(G130), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n630), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n818), .A2(new_n833), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n900), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n908), .B(new_n631), .ZN(new_n912));
  INV_X1    g487(.A(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(new_n899), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n898), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n898), .B1(new_n914), .B2(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n894), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n898), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n911), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n893), .A3(new_n915), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n882), .A2(new_n927), .A3(new_n573), .A4(new_n562), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n609), .B1(new_n929), .B2(new_n616), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n927), .B1(new_n620), .B2(new_n882), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT103), .B1(G299), .B2(new_n609), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n934), .A2(KEYINPUT41), .A3(new_n930), .A4(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(KEYINPUT105), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n878), .B(new_n625), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(new_n926), .C1(new_n931), .C2(new_n932), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n931), .B2(new_n932), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n934), .A2(KEYINPUT104), .A3(new_n930), .A4(new_n928), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n940), .B1(new_n945), .B2(new_n937), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(G303), .B(new_n751), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n950));
  NAND2_X1  g525(.A1(G288), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n514), .A2(G49), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n952), .A2(KEYINPUT106), .A3(new_n576), .A4(new_n577), .ZN(new_n953));
  AOI21_X1  g528(.A(G305), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n953), .A3(G305), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n949), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G303), .B(G290), .ZN(new_n958));
  INV_X1    g533(.A(new_n954), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n955), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT42), .Z(new_n962));
  AND2_X1   g537(.A1(new_n948), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n940), .B(KEYINPUT107), .C1(new_n945), .C2(new_n937), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n948), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n888), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(G868), .B2(new_n967), .ZN(G295));
  OAI21_X1  g543(.A(new_n966), .B1(G868), .B2(new_n967), .ZN(G331));
  NAND2_X1  g544(.A1(new_n526), .A2(new_n529), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT71), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G171), .B1(new_n973), .B2(new_n522), .ZN(new_n974));
  OAI211_X1 g549(.A(G171), .B(new_n522), .C1(new_n530), .C2(new_n531), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n974), .A2(new_n976), .B1(new_n876), .B2(new_n877), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n888), .A2(new_n547), .ZN(new_n979));
  NAND2_X1  g554(.A1(G286), .A2(G301), .ZN(new_n980));
  INV_X1    g555(.A(new_n877), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n975), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n878), .A2(KEYINPUT109), .A3(new_n980), .A4(new_n975), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n928), .A2(new_n930), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n934), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n961), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  OAI221_X1 g563(.A(KEYINPUT108), .B1(new_n876), .B2(new_n877), .C1(new_n974), .C2(new_n976), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n977), .A2(new_n990), .A3(new_n982), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n936), .A2(new_n939), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n992), .A3(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(new_n987), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G37), .B1(new_n999), .B2(new_n961), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT43), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n991), .A2(new_n989), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n944), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT41), .B1(new_n986), .B2(new_n934), .ZN(new_n1004));
  INV_X1    g579(.A(new_n935), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n984), .B(new_n983), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G37), .B1(new_n1007), .B2(new_n961), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n988), .A2(new_n992), .A3(KEYINPUT110), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT110), .B1(new_n988), .B2(new_n992), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1008), .B(KEYINPUT43), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n997), .B2(new_n1000), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1008), .B(new_n1015), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1019), .ZN(G397));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT112), .B(G40), .Z(new_n1023));
  OR3_X1    g598(.A1(new_n464), .A2(new_n467), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n493), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n485), .B2(new_n492), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT118), .A3(KEYINPUT45), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1027), .B2(new_n1025), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n464), .A2(new_n467), .A3(new_n1023), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1033), .A2(new_n789), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1022), .B1(new_n1040), .B2(G168), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1033), .A2(new_n789), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1034), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G286), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1021), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(G168), .A3(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(KEYINPUT51), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT62), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1040), .A2(G168), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT51), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1041), .A2(new_n1021), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1035), .A2(new_n1029), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n721), .A2(G1976), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1059), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n726), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G305), .A2(G1981), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1066), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1056), .A2(G8), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1063), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G166), .B2(new_n1022), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2090), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1027), .A2(new_n1025), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT111), .B(G1384), .Z(new_n1086));
  NAND3_X1  g661(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1035), .A3(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT113), .B(G1971), .Z(new_n1089));
  AOI22_X1  g664(.A1(new_n1039), .A2(new_n1084), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1083), .B1(new_n1022), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1039), .A2(new_n1084), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1022), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1076), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1098));
  INV_X1    g673(.A(G1961), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1088), .B2(G2078), .ZN(new_n1102));
  INV_X1    g677(.A(G2078), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT53), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1100), .B(new_n1102), .C1(new_n1033), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1097), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1050), .A2(new_n1055), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1076), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1066), .B(KEYINPUT117), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G288), .A2(G1976), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1113), .B2(new_n1073), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1040), .A2(new_n1022), .A3(G286), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1097), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(KEYINPUT63), .A3(new_n1076), .A4(new_n1116), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n620), .B2(KEYINPUT119), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  NAND3_X1  g701(.A1(G299), .A2(new_n1126), .A3(KEYINPUT57), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1085), .A2(new_n1035), .A3(new_n1087), .A4(new_n1128), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1125), .A2(new_n1131), .A3(new_n1129), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT121), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1123), .A2(new_n1137), .A3(new_n1127), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n772), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1056), .ZN(new_n1142));
  INV_X1    g717(.A(G2067), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n609), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1130), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT61), .B1(new_n1148), .B2(new_n1135), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT58), .B(G1341), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1088), .A2(G1996), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n548), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n609), .A2(KEYINPUT124), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1145), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1145), .A2(new_n1157), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n882), .B(KEYINPUT124), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1160), .A2(new_n1141), .A3(KEYINPUT60), .A4(new_n1144), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1150), .A2(new_n1155), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1125), .A2(new_n1129), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1130), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1147), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1105), .A2(G171), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT54), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1028), .A2(new_n1103), .A3(new_n1087), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1172), .A2(new_n1101), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1173));
  NAND2_X1  g748(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(KEYINPUT125), .B2(new_n1103), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(KEYINPUT125), .B2(new_n1103), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n468), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n493), .A2(new_n1086), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1025), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1179), .A3(new_n1087), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1173), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1171), .B1(new_n1181), .B2(G171), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1097), .B1(new_n1170), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1173), .A2(new_n1185), .A3(G301), .A4(new_n1180), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1100), .A2(G301), .A3(new_n1102), .A4(new_n1180), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT126), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1106), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1171), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1183), .A2(new_n1184), .A3(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1108), .B(new_n1121), .C1(new_n1169), .C2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1179), .A2(new_n1024), .ZN(new_n1193));
  INV_X1    g768(.A(new_n744), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n742), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1195), .A2(new_n748), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n802), .B(new_n1143), .ZN(new_n1197));
  INV_X1    g772(.A(G1996), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n833), .B(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n748), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(G290), .B(G1986), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1193), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1192), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT46), .Z(new_n1206));
  NAND3_X1  g781(.A1(new_n1197), .A2(new_n827), .A3(new_n832), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1206), .B1(new_n1207), .B2(new_n1193), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT47), .Z(new_n1209));
  NAND2_X1  g784(.A1(new_n1201), .A2(new_n1193), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1193), .A2(new_n754), .A3(new_n751), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT48), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1199), .A2(new_n1197), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1214), .A2(new_n1200), .B1(G2067), .B2(new_n802), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1193), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1209), .A2(new_n1213), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1204), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g793(.A(G319), .ZN(new_n1220));
  NOR2_X1   g794(.A1(G227), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1221), .B1(new_n713), .B2(new_n714), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n672), .B2(new_n673), .ZN(new_n1223));
  OAI211_X1 g797(.A(new_n924), .B(new_n1223), .C1(new_n1016), .C2(new_n1018), .ZN(G225));
  INV_X1    g798(.A(G225), .ZN(G308));
endmodule


