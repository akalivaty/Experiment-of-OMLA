

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n515) );
  NOR2_X1 U551 ( .A1(n742), .A2(n741), .ZN(n514) );
  XNOR2_X1 U552 ( .A(n710), .B(KEYINPUT30), .ZN(n711) );
  XNOR2_X1 U553 ( .A(n712), .B(n711), .ZN(n713) );
  OR2_X1 U554 ( .A1(n719), .A2(n718), .ZN(n731) );
  XNOR2_X1 U555 ( .A(n675), .B(KEYINPUT64), .ZN(n708) );
  OR2_X1 U556 ( .A1(n736), .A2(n735), .ZN(n789) );
  AND2_X1 U557 ( .A1(n789), .A2(n743), .ZN(n739) );
  AND2_X1 U558 ( .A1(n520), .A2(G2104), .ZN(n991) );
  NOR2_X1 U559 ( .A1(n643), .A2(G651), .ZN(n636) );
  XNOR2_X1 U560 ( .A(n516), .B(n515), .ZN(n519) );
  INV_X1 U561 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U562 ( .A1(G101), .A2(n991), .ZN(n516) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n517), .Z(n992) );
  NAND2_X1 U565 ( .A1(G137), .A2(n992), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n524) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n999) );
  NAND2_X1 U568 ( .A1(G113), .A2(n999), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n520), .ZN(n996) );
  NAND2_X1 U570 ( .A1(G125), .A2(n996), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n524), .A2(n523), .ZN(G160) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n627) );
  NAND2_X1 U574 ( .A1(G85), .A2(n627), .ZN(n526) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  INV_X1 U576 ( .A(G651), .ZN(n527) );
  NOR2_X1 U577 ( .A1(n643), .A2(n527), .ZN(n630) );
  NAND2_X1 U578 ( .A1(G72), .A2(n630), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U580 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n528), .Z(n641) );
  NAND2_X1 U582 ( .A1(G60), .A2(n641), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G47), .A2(n636), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  OR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(G290) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U587 ( .A1(n996), .A2(G123), .ZN(n534) );
  XNOR2_X1 U588 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n533) );
  XNOR2_X1 U589 ( .A(n534), .B(n533), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G99), .A2(n991), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G135), .A2(n992), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G111), .A2(n999), .ZN(n537) );
  XNOR2_X1 U594 ( .A(KEYINPUT77), .B(n537), .ZN(n538) );
  NOR2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n982) );
  XNOR2_X1 U597 ( .A(G2096), .B(n982), .ZN(n542) );
  OR2_X1 U598 ( .A1(G2100), .A2(n542), .ZN(G156) );
  INV_X1 U599 ( .A(G108), .ZN(G238) );
  INV_X1 U600 ( .A(G120), .ZN(G236) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(n627), .A2(G90), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n543), .B(KEYINPUT68), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G77), .A2(n630), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(KEYINPUT9), .B(n546), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n641), .A2(G64), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n547), .B(KEYINPUT66), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G52), .A2(n636), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT67), .B(n550), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(G301) );
  INV_X1 U614 ( .A(G301), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n627), .A2(G89), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U617 ( .A1(G76), .A2(n630), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G63), .A2(n641), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G51), .A2(n636), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U626 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U627 ( .A1(n991), .A2(G102), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT86), .ZN(n565) );
  NAND2_X1 U629 ( .A1(G126), .A2(n996), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G138), .A2(n992), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G114), .A2(n999), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(G164) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G567), .ZN(n669) );
  NOR2_X1 U638 ( .A1(n669), .A2(G223), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n571), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U640 ( .A1(n641), .A2(G56), .ZN(n572) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n572), .Z(n578) );
  NAND2_X1 U642 ( .A1(n627), .A2(G81), .ZN(n573) );
  XNOR2_X1 U643 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G68), .A2(n630), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U648 ( .A(KEYINPUT70), .B(n579), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n636), .A2(G43), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT71), .B(n580), .Z(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n1009) );
  INV_X1 U652 ( .A(G860), .ZN(n604) );
  OR2_X1 U653 ( .A1(n1009), .A2(n604), .ZN(G153) );
  NAND2_X1 U654 ( .A1(G301), .A2(G868), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT72), .ZN(n594) );
  NAND2_X1 U656 ( .A1(G92), .A2(n627), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G66), .A2(n641), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT73), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G79), .A2(n630), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n636), .A2(G54), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT74), .B(n589), .Z(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT15), .B(n592), .Z(n1010) );
  OR2_X1 U666 ( .A1(G868), .A2(n1010), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U668 ( .A1(G65), .A2(n641), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G53), .A2(n636), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G91), .A2(n627), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G78), .A2(n630), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n849) );
  INV_X1 U675 ( .A(G868), .ZN(n653) );
  NAND2_X1 U676 ( .A1(n849), .A2(n653), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT75), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n653), .A2(G286), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n604), .A2(G559), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n605), .A2(n1010), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n1009), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G868), .A2(n1010), .ZN(n607) );
  NOR2_X1 U685 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G282) );
  XNOR2_X1 U687 ( .A(n1009), .B(KEYINPUT78), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n1010), .A2(G559), .ZN(n610) );
  XNOR2_X1 U689 ( .A(n611), .B(n610), .ZN(n651) );
  NOR2_X1 U690 ( .A1(n651), .A2(G860), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G93), .A2(n627), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G80), .A2(n630), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G55), .A2(n636), .ZN(n614) );
  XNOR2_X1 U695 ( .A(KEYINPUT79), .B(n614), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n641), .A2(G67), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n654) );
  XOR2_X1 U699 ( .A(n654), .B(KEYINPUT80), .Z(n619) );
  XNOR2_X1 U700 ( .A(n620), .B(n619), .ZN(G145) );
  NAND2_X1 U701 ( .A1(G88), .A2(n627), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G75), .A2(n630), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G62), .A2(n641), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G50), .A2(n636), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(G166) );
  NAND2_X1 U708 ( .A1(G86), .A2(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G61), .A2(n641), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n630), .A2(G73), .ZN(n631) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(G48), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G49), .A2(n636), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT81), .B(n639), .Z(n640) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT82), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n643), .A2(G87), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(G288) );
  XNOR2_X1 U724 ( .A(G290), .B(KEYINPUT19), .ZN(n647) );
  XNOR2_X1 U725 ( .A(G166), .B(n849), .ZN(n646) );
  XNOR2_X1 U726 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(G305), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(n654), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n650), .B(G288), .ZN(n1013) );
  XOR2_X1 U730 ( .A(n1013), .B(n651), .Z(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n656) );
  NOR2_X1 U732 ( .A1(G868), .A2(n654), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n660), .A2(G2072), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT83), .B(n661), .Z(G158) );
  XNOR2_X1 U740 ( .A(KEYINPUT84), .B(G44), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n662), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U742 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n663) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n663), .Z(n664) );
  NOR2_X1 U745 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G96), .A2(n665), .ZN(n957) );
  NAND2_X1 U747 ( .A1(G2106), .A2(n957), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(KEYINPUT85), .ZN(n671) );
  NOR2_X1 U749 ( .A1(G236), .A2(G238), .ZN(n667) );
  NAND2_X1 U750 ( .A1(G69), .A2(n667), .ZN(n668) );
  NOR2_X1 U751 ( .A1(G237), .A2(n668), .ZN(n959) );
  NOR2_X1 U752 ( .A1(n669), .A2(n959), .ZN(n670) );
  NOR2_X1 U753 ( .A1(n671), .A2(n670), .ZN(G319) );
  INV_X1 U754 ( .A(G319), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U756 ( .A1(n673), .A2(n672), .ZN(n840) );
  NAND2_X1 U757 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  AND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n674) );
  NOR2_X1 U760 ( .A1(G164), .A2(G1384), .ZN(n773) );
  NAND2_X1 U761 ( .A1(n674), .A2(n773), .ZN(n675) );
  INV_X1 U762 ( .A(n708), .ZN(n701) );
  NAND2_X1 U763 ( .A1(G2072), .A2(n701), .ZN(n676) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(n676), .Z(n678) );
  INV_X1 U765 ( .A(n701), .ZN(n721) );
  NAND2_X1 U766 ( .A1(n721), .A2(G1956), .ZN(n677) );
  NAND2_X1 U767 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U768 ( .A(KEYINPUT92), .B(n679), .Z(n694) );
  NOR2_X1 U769 ( .A1(n849), .A2(n694), .ZN(n681) );
  XNOR2_X1 U770 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n680) );
  XNOR2_X1 U771 ( .A(n681), .B(n680), .ZN(n698) );
  NAND2_X1 U772 ( .A1(G1996), .A2(n701), .ZN(n682) );
  XNOR2_X1 U773 ( .A(n682), .B(KEYINPUT26), .ZN(n684) );
  NAND2_X1 U774 ( .A1(G1341), .A2(n708), .ZN(n683) );
  NAND2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U776 ( .A(KEYINPUT94), .B(n685), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n686), .A2(n1009), .ZN(n691) );
  NAND2_X1 U778 ( .A1(n691), .A2(n1010), .ZN(n690) );
  NOR2_X1 U779 ( .A1(n721), .A2(G2067), .ZN(n688) );
  NOR2_X1 U780 ( .A1(G1348), .A2(n701), .ZN(n687) );
  NOR2_X1 U781 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n693) );
  OR2_X1 U783 ( .A1(n1010), .A2(n691), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n849), .A2(n694), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U788 ( .A(n699), .B(KEYINPUT29), .ZN(n706) );
  XOR2_X1 U789 ( .A(G2078), .B(KEYINPUT25), .Z(n700) );
  XNOR2_X1 U790 ( .A(KEYINPUT90), .B(n700), .ZN(n889) );
  NAND2_X1 U791 ( .A1(n701), .A2(n889), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n721), .A2(G1961), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U794 ( .A(KEYINPUT91), .B(n704), .ZN(n707) );
  AND2_X1 U795 ( .A1(G171), .A2(n707), .ZN(n705) );
  NOR2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n719) );
  NOR2_X1 U797 ( .A1(G171), .A2(n707), .ZN(n715) );
  NAND2_X1 U798 ( .A1(n708), .A2(G8), .ZN(n797) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n797), .ZN(n734) );
  NOR2_X1 U800 ( .A1(n721), .A2(G2084), .ZN(n732) );
  NOR2_X1 U801 ( .A1(n734), .A2(n732), .ZN(n709) );
  NAND2_X1 U802 ( .A1(G8), .A2(n709), .ZN(n712) );
  INV_X1 U803 ( .A(KEYINPUT95), .ZN(n710) );
  NOR2_X1 U804 ( .A1(G168), .A2(n713), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT96), .B(n716), .ZN(n717) );
  XNOR2_X1 U807 ( .A(KEYINPUT31), .B(n717), .ZN(n718) );
  AND2_X1 U808 ( .A1(G286), .A2(G8), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n731), .A2(n720), .ZN(n728) );
  INV_X1 U810 ( .A(G8), .ZN(n726) );
  NOR2_X1 U811 ( .A1(n721), .A2(G2090), .ZN(n723) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n797), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n724), .A2(G303), .ZN(n725) );
  OR2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U817 ( .A(n729), .B(KEYINPUT98), .ZN(n730) );
  XNOR2_X1 U818 ( .A(KEYINPUT32), .B(n730), .ZN(n788) );
  XNOR2_X1 U819 ( .A(n731), .B(KEYINPUT97), .ZN(n736) );
  AND2_X1 U820 ( .A1(n732), .A2(G8), .ZN(n733) );
  OR2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n735) );
  INV_X1 U822 ( .A(KEYINPUT33), .ZN(n738) );
  NAND2_X1 U823 ( .A1(G288), .A2(G1976), .ZN(n737) );
  XOR2_X1 U824 ( .A(KEYINPUT101), .B(n737), .Z(n922) );
  AND2_X1 U825 ( .A1(n738), .A2(n922), .ZN(n743) );
  NAND2_X1 U826 ( .A1(n788), .A2(n739), .ZN(n753) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n910) );
  INV_X1 U828 ( .A(n797), .ZN(n741) );
  NAND2_X1 U829 ( .A1(n910), .A2(n741), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n740), .A2(KEYINPUT33), .ZN(n749) );
  INV_X1 U831 ( .A(n749), .ZN(n742) );
  INV_X1 U832 ( .A(n743), .ZN(n748) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n744) );
  XOR2_X1 U834 ( .A(n744), .B(KEYINPUT99), .Z(n745) );
  NOR2_X1 U835 ( .A1(n910), .A2(n745), .ZN(n746) );
  XNOR2_X1 U836 ( .A(n746), .B(KEYINPUT100), .ZN(n747) );
  OR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n750) );
  AND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  OR2_X1 U839 ( .A1(n514), .A2(n751), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U841 ( .A(n754), .B(KEYINPUT102), .ZN(n787) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n906) );
  XNOR2_X1 U843 ( .A(KEYINPUT87), .B(G1986), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(G290), .ZN(n918) );
  NAND2_X1 U845 ( .A1(n996), .A2(G119), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G131), .A2(n992), .ZN(n756) );
  XOR2_X1 U847 ( .A(KEYINPUT89), .B(n756), .Z(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G95), .A2(n991), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G107), .A2(n999), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n980) );
  INV_X1 U853 ( .A(G1991), .ZN(n803) );
  NOR2_X1 U854 ( .A1(n980), .A2(n803), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n991), .A2(G105), .ZN(n763) );
  XNOR2_X1 U856 ( .A(n763), .B(KEYINPUT38), .ZN(n765) );
  NAND2_X1 U857 ( .A1(G129), .A2(n996), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G141), .A2(n992), .ZN(n767) );
  NAND2_X1 U860 ( .A1(G117), .A2(n999), .ZN(n766) );
  NAND2_X1 U861 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U862 ( .A1(n769), .A2(n768), .ZN(n984) );
  INV_X1 U863 ( .A(G1996), .ZN(n802) );
  NOR2_X1 U864 ( .A1(n984), .A2(n802), .ZN(n770) );
  NOR2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n865) );
  NAND2_X1 U866 ( .A1(n918), .A2(n865), .ZN(n774) );
  NAND2_X1 U867 ( .A1(G160), .A2(G40), .ZN(n772) );
  NOR2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n817) );
  NAND2_X1 U869 ( .A1(n774), .A2(n817), .ZN(n785) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n813) );
  NAND2_X1 U871 ( .A1(G116), .A2(n999), .ZN(n776) );
  NAND2_X1 U872 ( .A1(G128), .A2(n996), .ZN(n775) );
  NAND2_X1 U873 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U874 ( .A(n777), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U875 ( .A1(G104), .A2(n991), .ZN(n779) );
  NAND2_X1 U876 ( .A1(G140), .A2(n992), .ZN(n778) );
  NAND2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U878 ( .A(KEYINPUT34), .B(n780), .Z(n781) );
  NAND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U880 ( .A(n783), .B(KEYINPUT36), .Z(n1005) );
  OR2_X1 U881 ( .A1(n813), .A2(n1005), .ZN(n784) );
  XOR2_X1 U882 ( .A(KEYINPUT88), .B(n784), .Z(n867) );
  NAND2_X1 U883 ( .A1(n817), .A2(n867), .ZN(n811) );
  AND2_X1 U884 ( .A1(n785), .A2(n811), .ZN(n799) );
  AND2_X1 U885 ( .A1(n906), .A2(n799), .ZN(n786) );
  AND2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n822) );
  NAND2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n792) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n790) );
  NAND2_X1 U889 ( .A1(G8), .A2(n790), .ZN(n791) );
  NAND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n794) );
  AND2_X1 U891 ( .A1(n797), .A2(n799), .ZN(n793) );
  AND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n801) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U894 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  NOR2_X1 U895 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n820) );
  AND2_X1 U898 ( .A1(n802), .A2(n984), .ZN(n872) );
  INV_X1 U899 ( .A(n865), .ZN(n808) );
  AND2_X1 U900 ( .A1(n980), .A2(n803), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT104), .ZN(n863) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n805) );
  XOR2_X1 U903 ( .A(n805), .B(KEYINPUT103), .Z(n806) );
  NOR2_X1 U904 ( .A1(n863), .A2(n806), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n872), .A2(n809), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n1005), .A2(n813), .ZN(n869) );
  NAND2_X1 U910 ( .A1(n814), .A2(n869), .ZN(n815) );
  XOR2_X1 U911 ( .A(KEYINPUT105), .B(n815), .Z(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U913 ( .A(KEYINPUT106), .B(n818), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U916 ( .A(n823), .B(KEYINPUT40), .Z(G329) );
  XOR2_X1 U917 ( .A(G2454), .B(G2427), .Z(n825) );
  XNOR2_X1 U918 ( .A(KEYINPUT108), .B(KEYINPUT107), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n825), .B(n824), .ZN(n835) );
  XOR2_X1 U920 ( .A(G2443), .B(G2446), .Z(n827) );
  XNOR2_X1 U921 ( .A(G1348), .B(G2438), .ZN(n826) );
  XNOR2_X1 U922 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U923 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n829) );
  XNOR2_X1 U924 ( .A(G2430), .B(G2435), .ZN(n828) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U926 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U927 ( .A(G1341), .B(G2451), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n836), .A2(G14), .ZN(n1017) );
  XNOR2_X1 U931 ( .A(KEYINPUT111), .B(n1017), .ZN(G401) );
  INV_X1 U932 ( .A(G223), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U935 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G188) );
  NAND2_X1 U939 ( .A1(G100), .A2(n991), .ZN(n842) );
  NAND2_X1 U940 ( .A1(G112), .A2(n999), .ZN(n841) );
  NAND2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n848) );
  NAND2_X1 U942 ( .A1(n996), .A2(G124), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n843), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U944 ( .A1(G136), .A2(n992), .ZN(n844) );
  NAND2_X1 U945 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(KEYINPUT115), .B(n846), .Z(n847) );
  NOR2_X1 U947 ( .A1(n848), .A2(n847), .ZN(G162) );
  INV_X1 U948 ( .A(n849), .ZN(G299) );
  INV_X1 U949 ( .A(KEYINPUT55), .ZN(n901) );
  NAND2_X1 U950 ( .A1(G103), .A2(n991), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G139), .A2(n992), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n851), .A2(n850), .ZN(n857) );
  NAND2_X1 U953 ( .A1(n996), .A2(G127), .ZN(n852) );
  XOR2_X1 U954 ( .A(KEYINPUT117), .B(n852), .Z(n854) );
  NAND2_X1 U955 ( .A1(n999), .A2(G115), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(KEYINPUT47), .B(n855), .Z(n856) );
  NOR2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n981) );
  XOR2_X1 U959 ( .A(G2072), .B(n981), .Z(n859) );
  XOR2_X1 U960 ( .A(G164), .B(G2078), .Z(n858) );
  NOR2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(KEYINPUT50), .B(n860), .Z(n878) );
  XNOR2_X1 U963 ( .A(G160), .B(G2084), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n861), .A2(n982), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT120), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n875) );
  XOR2_X1 U970 ( .A(G2090), .B(G162), .Z(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT51), .ZN(n874) );
  NOR2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT121), .B(n876), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n879), .B(KEYINPUT122), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n880), .B(KEYINPUT52), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n901), .A2(n881), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n882), .A2(G29), .ZN(n931) );
  XNOR2_X1 U980 ( .A(G2084), .B(G34), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(KEYINPUT54), .ZN(n885) );
  XNOR2_X1 U982 ( .A(G35), .B(G2090), .ZN(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n899) );
  XOR2_X1 U984 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n897) );
  XOR2_X1 U985 ( .A(G2067), .B(G26), .Z(n886) );
  NAND2_X1 U986 ( .A1(n886), .A2(G28), .ZN(n895) );
  XNOR2_X1 U987 ( .A(G2072), .B(G33), .ZN(n888) );
  XNOR2_X1 U988 ( .A(G25), .B(G1991), .ZN(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n889), .B(G27), .ZN(n891) );
  XNOR2_X1 U991 ( .A(G1996), .B(G32), .ZN(n890) );
  NOR2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  NOR2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n898) );
  NAND2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  INV_X1 U998 ( .A(G29), .ZN(n902) );
  NAND2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G11), .A2(n904), .ZN(n929) );
  XOR2_X1 U1001 ( .A(KEYINPUT56), .B(G16), .Z(n927) );
  XNOR2_X1 U1002 ( .A(G168), .B(G1966), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(KEYINPUT124), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(KEYINPUT57), .ZN(n912) );
  XOR2_X1 U1006 ( .A(G1961), .B(G171), .Z(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n925) );
  XNOR2_X1 U1009 ( .A(G303), .B(G1971), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(G299), .B(G1956), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(G1341), .B(KEYINPUT125), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n915), .B(n1009), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G1348), .B(n1010), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1022 ( .A1(n931), .A2(n930), .ZN(n955) );
  XOR2_X1 U1023 ( .A(G1986), .B(G24), .Z(n935) );
  XNOR2_X1 U1024 ( .A(G1971), .B(G22), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(G23), .B(G1976), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(KEYINPUT58), .B(n936), .ZN(n951) );
  XOR2_X1 U1029 ( .A(G1961), .B(G5), .Z(n949) );
  XNOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(n937), .B(G4), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(G20), .B(G1956), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT60), .B(n944), .Z(n946) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G21), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT126), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1044 ( .A(KEYINPUT61), .B(n952), .Z(n953) );
  NOR2_X1 U1045 ( .A1(G16), .A2(n953), .ZN(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1049 ( .A(G96), .ZN(G221) );
  INV_X1 U1050 ( .A(n957), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(G261) );
  INV_X1 U1052 ( .A(G261), .ZN(G325) );
  XOR2_X1 U1053 ( .A(KEYINPUT113), .B(G2474), .Z(n961) );
  XNOR2_X1 U1054 ( .A(G1961), .B(G1976), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(n962), .B(KEYINPUT41), .Z(n964) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G1991), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT114), .B(G1986), .Z(n966) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G1956), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1062 ( .A(n968), .B(n967), .Z(n970) );
  XNOR2_X1 U1063 ( .A(G1996), .B(G1981), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n970), .B(n969), .ZN(G229) );
  XOR2_X1 U1065 ( .A(G2100), .B(G2096), .Z(n972) );
  XNOR2_X1 U1066 ( .A(G2090), .B(KEYINPUT112), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1068 ( .A(n973), .B(KEYINPUT42), .Z(n975) );
  XNOR2_X1 U1069 ( .A(G2072), .B(KEYINPUT43), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n975), .B(n974), .ZN(n979) );
  XOR2_X1 U1071 ( .A(G2678), .B(G2067), .Z(n977) );
  XNOR2_X1 U1072 ( .A(G2084), .B(G2078), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n979), .B(n978), .ZN(G227) );
  XOR2_X1 U1075 ( .A(n981), .B(n980), .Z(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(n982), .ZN(n988) );
  XOR2_X1 U1077 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n986) );
  XNOR2_X1 U1078 ( .A(n984), .B(KEYINPUT118), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1080 ( .A(n988), .B(n987), .Z(n990) );
  XNOR2_X1 U1081 ( .A(G160), .B(G164), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n990), .B(n989), .ZN(n1004) );
  NAND2_X1 U1083 ( .A1(G106), .A2(n991), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(G142), .A2(n992), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT45), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(G130), .A2(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n999), .A2(G118), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT116), .B(n1000), .Z(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(n1004), .B(n1003), .Z(n1007) );
  XOR2_X1 U1093 ( .A(n1005), .B(G162), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(n1007), .B(n1006), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(G37), .A2(n1008), .ZN(G395) );
  XNOR2_X1 U1096 ( .A(n1009), .B(KEYINPUT119), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G171), .B(n1010), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1012), .B(n1011), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(G286), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1100 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(G37), .A2(n1016), .ZN(G397) );
  NAND2_X1 U1102 ( .A1(G319), .A2(n1017), .ZN(n1020) );
  NOR2_X1 U1103 ( .A1(G229), .A2(G227), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT49), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(G395), .A2(G397), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(G225) );
  INV_X1 U1108 ( .A(G225), .ZN(G308) );
  INV_X1 U1109 ( .A(G69), .ZN(G235) );
endmodule

