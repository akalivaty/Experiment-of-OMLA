//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G113), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n191), .B(new_n193), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n193), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT2), .B(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n200), .A3(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G104), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(G107), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n206), .A2(KEYINPUT3), .A3(G107), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(G107), .B1(new_n207), .B2(new_n209), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n210), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G101), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT4), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n205), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n215), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n223), .B1(new_n215), .B2(new_n226), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n189), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n218), .A2(new_n220), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n208), .A2(G104), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n232), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n206), .B2(G107), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n213), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT82), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n219), .B1(new_n213), .B2(new_n232), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n231), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n190), .A3(G116), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n250));
  OAI21_X1  g064(.A(G113), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n250), .B2(new_n249), .ZN(new_n252));
  INV_X1    g066(.A(new_n198), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n247), .A2(new_n197), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n215), .A2(new_n226), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT80), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n215), .A2(new_n223), .A3(new_n226), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n211), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g075(.A(new_n220), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n216), .A3(KEYINPUT4), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n260), .A2(KEYINPUT86), .A3(new_n205), .A4(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n230), .A2(new_n256), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G122), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT88), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n188), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n230), .A2(new_n256), .A3(new_n265), .A4(new_n267), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT89), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT90), .ZN(new_n275));
  INV_X1    g089(.A(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT1), .B1(new_n278), .B2(G146), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(G128), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n277), .B(new_n279), .C1(KEYINPUT1), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n277), .A2(new_n279), .A3(new_n289), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n280), .A2(new_n291), .A3(KEYINPUT64), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n288), .B1(new_n287), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G224), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G953), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT91), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n298), .B(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n266), .A2(new_n188), .A3(new_n268), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n305), .B(new_n269), .C1(new_n272), .C2(new_n273), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n275), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n273), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n270), .A2(new_n271), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT7), .B1(new_n299), .B2(G953), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n298), .B(new_n310), .Z(new_n311));
  NOR3_X1   g125(.A1(new_n237), .A2(new_n240), .A3(KEYINPUT82), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n245), .B1(new_n242), .B2(new_n244), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n263), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n255), .A2(new_n197), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT94), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT92), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n254), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n253), .A2(KEYINPUT92), .A3(KEYINPUT5), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n252), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n197), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT93), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(KEYINPUT93), .A3(new_n197), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n247), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n327), .A3(new_n315), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n267), .B(KEYINPUT8), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n311), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n308), .A2(new_n309), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G210), .B1(G237), .B2(G902), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n307), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n307), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n187), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G469), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G140), .ZN(new_n341));
  INV_X1    g155(.A(G953), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(G227), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G134), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT65), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G137), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT11), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n346), .A2(new_n348), .A3(G137), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT66), .A2(G137), .ZN(new_n355));
  AND2_X1   g169(.A1(KEYINPUT11), .A2(G134), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G131), .B1(new_n351), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT11), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT65), .B(G134), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(G137), .ZN(new_n362));
  INV_X1    g176(.A(G131), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n352), .A4(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT70), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n359), .A2(KEYINPUT70), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n286), .B(new_n263), .C1(new_n312), .C2(new_n313), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n241), .A2(new_n246), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n286), .B1(new_n372), .B2(new_n263), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT12), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n314), .A2(new_n285), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n370), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n359), .B2(new_n364), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n374), .A2(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n296), .A2(new_n295), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT64), .B1(new_n280), .B2(new_n291), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n294), .A2(KEYINPUT69), .A3(new_n295), .A4(new_n296), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n260), .A3(new_n264), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n370), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n359), .A2(KEYINPUT70), .A3(new_n364), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT70), .B1(new_n359), .B2(new_n364), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n286), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n387), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n344), .B1(new_n380), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n344), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT84), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(KEYINPUT84), .A3(new_n397), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n387), .A2(new_n389), .A3(new_n393), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n369), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n396), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G902), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n340), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT85), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n407));
  INV_X1    g221(.A(new_n398), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n401), .A3(new_n399), .ZN(new_n409));
  AOI21_X1  g223(.A(G902), .B1(new_n409), .B2(new_n396), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(new_n340), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n394), .A2(new_n397), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n380), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n397), .B1(new_n401), .B2(new_n394), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n340), .B(new_n404), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n406), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT9), .B(G234), .ZN(new_n417));
  OAI21_X1  g231(.A(G221), .B1(new_n417), .B2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G125), .B(G140), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g235(.A(G140), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G125), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(KEYINPUT16), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n276), .ZN(new_n425));
  NOR2_X1   g239(.A1(G237), .A2(G953), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n426), .A2(G143), .A3(G214), .ZN(new_n427));
  AOI21_X1  g241(.A(G143), .B1(new_n426), .B2(G214), .ZN(new_n428));
  OAI21_X1  g242(.A(G131), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(G214), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n278), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n426), .A2(G143), .A3(G214), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n363), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n421), .B(G146), .C1(KEYINPUT16), .C2(new_n423), .ZN(new_n436));
  OAI211_X1 g250(.A(KEYINPUT17), .B(G131), .C1(new_n427), .C2(new_n428), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n425), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n206), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n420), .A2(KEYINPUT75), .A3(new_n276), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT75), .B1(new_n420), .B2(new_n276), .ZN(new_n442));
  OAI22_X1  g256(.A1(new_n441), .A2(new_n442), .B1(new_n276), .B2(new_n420), .ZN(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n431), .A2(new_n432), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT18), .B(G131), .C1(new_n427), .C2(new_n428), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n438), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n420), .A2(KEYINPUT19), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n420), .A2(KEYINPUT19), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n276), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n429), .A2(new_n433), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n436), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n440), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT96), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(G475), .A2(G902), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n447), .A2(new_n453), .ZN(new_n457));
  INV_X1    g271(.A(new_n440), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n438), .A2(new_n440), .A3(new_n447), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n461), .ZN(new_n465));
  NOR3_X1   g279(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT98), .ZN(new_n469));
  INV_X1    g283(.A(G475), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n440), .B1(new_n438), .B2(new_n447), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n448), .A2(new_n471), .A3(KEYINPUT97), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n471), .B2(KEYINPUT97), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n468), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n463), .A2(KEYINPUT20), .B1(new_n465), .B2(new_n466), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT98), .B1(new_n477), .B2(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(G116), .B(G122), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(G107), .B(new_n480), .C1(new_n482), .C2(KEYINPUT14), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n233), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n278), .A2(G128), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n283), .A2(G143), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n361), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n361), .B1(new_n485), .B2(new_n486), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n483), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n481), .B(new_n233), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n485), .A2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(G134), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n496), .A3(new_n487), .ZN(new_n497));
  INV_X1    g311(.A(G217), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n417), .A2(new_n498), .A3(G953), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n490), .B2(new_n497), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n404), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT99), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(KEYINPUT99), .B(new_n404), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(G478), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n505), .A2(new_n506), .A3(G478), .ZN(new_n508));
  OR3_X1    g322(.A1(new_n507), .A2(KEYINPUT100), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT100), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(G234), .A2(G237), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n512), .A2(G952), .A3(new_n342), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT21), .B(G898), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT101), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n512), .A2(G902), .A3(G953), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n479), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n339), .A2(new_n419), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G234), .ZN(new_n522));
  OAI21_X1  g336(.A(G217), .B1(new_n522), .B2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n425), .A2(new_n436), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n190), .A2(G128), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n283), .A2(KEYINPUT23), .A3(G119), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n190), .A2(G128), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(KEYINPUT23), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n283), .A2(G119), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n529), .A2(G110), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n529), .A2(G110), .B1(new_n531), .B2(new_n533), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(new_n436), .C1(new_n442), .C2(new_n441), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n342), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT76), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n538), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n524), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n549), .B2(new_n548), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n523), .A2(new_n404), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT67), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n382), .A2(new_n383), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n349), .A2(new_n350), .ZN(new_n558));
  INV_X1    g372(.A(new_n355), .ZN(new_n559));
  NOR2_X1   g373(.A1(KEYINPUT66), .A2(G137), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n345), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n363), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n285), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n365), .A2(new_n557), .B1(new_n563), .B2(new_n364), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n556), .B1(new_n564), .B2(KEYINPUT30), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n297), .B1(new_n364), .B2(new_n359), .ZN(new_n567));
  INV_X1    g381(.A(new_n562), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n568), .A2(new_n364), .A3(new_n286), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT67), .B(new_n566), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n569), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n384), .A2(new_n385), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT30), .B(new_n572), .C1(new_n392), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n205), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n572), .B(new_n204), .C1(new_n392), .C2(new_n573), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n369), .A2(new_n386), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n579), .A2(KEYINPUT71), .A3(new_n572), .A4(new_n204), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n426), .A2(G210), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT27), .Z(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT26), .B(G101), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n582), .B(new_n583), .Z(new_n584));
  NAND4_X1  g398(.A1(new_n575), .A2(new_n578), .A3(new_n580), .A4(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT72), .B1(new_n585), .B2(KEYINPUT31), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(KEYINPUT31), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n205), .B1(new_n567), .B2(new_n569), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n578), .A2(new_n590), .A3(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT28), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n569), .B1(new_n369), .B2(new_n386), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT28), .B1(new_n593), .B2(new_n204), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n584), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT73), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n591), .B2(KEYINPUT28), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT73), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n599), .A2(new_n600), .A3(new_n584), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n588), .B(new_n589), .C1(new_n598), .C2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(G472), .A2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT32), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n603), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n605), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT29), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n597), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n609), .B(new_n611), .C1(new_n596), .C2(new_n597), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n578), .B(new_n580), .C1(new_n204), .C2(new_n593), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n594), .B1(new_n613), .B2(KEYINPUT28), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n597), .A2(new_n609), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n602), .A2(new_n608), .B1(new_n617), .B2(G472), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n555), .B1(new_n606), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n521), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  NOR2_X1   g435(.A1(new_n500), .A2(new_n501), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n490), .A2(new_n497), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(KEYINPUT102), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n622), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G478), .ZN(new_n627));
  INV_X1    g441(.A(G478), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n404), .ZN(new_n629));
  INV_X1    g443(.A(new_n502), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n628), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n476), .B2(new_n478), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n339), .A2(new_n518), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n416), .A2(new_n418), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n602), .B2(new_n404), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n588), .A2(new_n589), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n596), .A2(KEYINPUT73), .A3(new_n597), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n600), .B1(new_n599), .B2(new_n584), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n607), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n638), .A2(new_n643), .A3(new_n555), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n635), .A2(new_n636), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n602), .A2(new_n404), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  INV_X1    g463(.A(new_n555), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n636), .A2(new_n649), .A3(new_n604), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n187), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n307), .A2(new_n335), .ZN(new_n653));
  INV_X1    g467(.A(new_n336), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n307), .A2(new_n335), .A3(new_n336), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n518), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n474), .B1(new_n659), .B2(new_n464), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n511), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT35), .B(G107), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n543), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n538), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n553), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n551), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(G902), .B1(new_n639), .B2(new_n642), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n604), .B(new_n670), .C1(new_n671), .C2(new_n637), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n649), .A2(KEYINPUT103), .A3(new_n604), .A4(new_n670), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n521), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n513), .B1(new_n517), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n679), .B1(new_n661), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n681), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n511), .A2(KEYINPUT104), .A3(new_n660), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n670), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n606), .B2(new_n618), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n339), .A2(new_n419), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XOR2_X1   g503(.A(new_n681), .B(KEYINPUT39), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n636), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n602), .A2(new_n608), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n610), .A2(new_n584), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n695), .B(new_n404), .C1(new_n584), .C2(new_n613), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n694), .B(new_n697), .C1(new_n643), .C2(KEYINPUT32), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n479), .A2(new_n511), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n337), .A2(new_n338), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT38), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT38), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n337), .B2(new_n338), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n670), .A2(new_n652), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n693), .A2(new_n701), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  NAND2_X1  g524(.A1(new_n606), .A2(new_n618), .ZN(new_n711));
  INV_X1    g525(.A(new_n632), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n479), .A2(new_n712), .A3(new_n683), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n687), .A2(new_n711), .A3(new_n670), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  OAI21_X1  g530(.A(new_n404), .B1(new_n413), .B2(new_n414), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G469), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n418), .A3(new_n415), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n635), .A2(new_n619), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT41), .B(G113), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G15));
  NOR2_X1   g538(.A1(new_n339), .A2(new_n518), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n619), .A2(new_n725), .A3(new_n662), .A4(new_n720), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  AOI211_X1 g541(.A(new_n652), .B(new_n719), .C1(new_n655), .C2(new_n656), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n711), .A3(new_n519), .A4(new_n670), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  XOR2_X1   g544(.A(new_n585), .B(KEYINPUT31), .Z(new_n731));
  OR2_X1    g545(.A1(new_n614), .A2(new_n584), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n607), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n638), .A2(new_n555), .A3(new_n733), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n652), .B(new_n699), .C1(new_n655), .C2(new_n656), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n719), .A2(new_n518), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT106), .B(G122), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G24));
  INV_X1    g553(.A(new_n670), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n638), .A2(new_n740), .A3(new_n733), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n633), .A2(new_n742), .A3(new_n683), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n742), .B1(new_n633), .B2(new_n683), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(new_n728), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NAND3_X1  g561(.A1(new_n655), .A2(new_n187), .A3(new_n656), .ZN(new_n748));
  INV_X1    g562(.A(new_n415), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n418), .B1(new_n405), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n752), .B(new_n418), .C1(new_n405), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n619), .A2(new_n755), .A3(new_n745), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT32), .B1(new_n602), .B2(new_n603), .ZN(new_n759));
  INV_X1    g573(.A(new_n608), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n639), .B2(new_n642), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n763), .B(new_n694), .C1(new_n643), .C2(KEYINPUT32), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n617), .A2(G472), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n633), .A2(new_n742), .A3(new_n683), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT42), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n748), .A2(new_n754), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n650), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n758), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  NAND2_X1  g587(.A1(new_n682), .A2(new_n684), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n619), .A2(new_n755), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n780));
  OAI22_X1  g594(.A1(new_n479), .A2(new_n632), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n476), .A2(new_n478), .A3(new_n712), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n780), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n649), .A2(new_n604), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n786), .A3(new_n670), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n748), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n340), .B1(new_n403), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n409), .A2(KEYINPUT45), .A3(new_n396), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n791), .A2(new_n792), .B1(G469), .B2(G902), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(KEYINPUT46), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n415), .B1(new_n793), .B2(KEYINPUT46), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n418), .B(new_n690), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n786), .A4(new_n670), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n789), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(G137), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G39));
  OAI21_X1  g615(.A(new_n418), .B1(new_n794), .B2(new_n795), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT47), .B(new_n418), .C1(new_n794), .C2(new_n795), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n337), .A2(new_n338), .A3(new_n652), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n711), .A2(new_n650), .A3(new_n713), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NOR2_X1   g624(.A1(G952), .A2(G953), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT121), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n718), .A2(new_n415), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n804), .B(new_n805), .C1(new_n418), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n783), .A2(new_n513), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n734), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n748), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n807), .A2(KEYINPUT117), .A3(new_n720), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n748), .B2(new_n719), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n513), .A3(new_n741), .A4(new_n783), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n698), .A2(new_n555), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n479), .A2(new_n712), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n513), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n719), .A2(new_n187), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n703), .B2(new_n705), .ZN(new_n830));
  AND4_X1   g644(.A1(KEYINPUT50), .A2(new_n830), .A3(new_n734), .A4(new_n815), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n734), .A2(new_n815), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT50), .B1(new_n832), .B2(new_n830), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n824), .B(new_n827), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n819), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n833), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n830), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n824), .A4(new_n827), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT51), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n823), .A2(new_n513), .A3(new_n783), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n766), .A2(new_n650), .ZN(new_n843));
  NOR2_X1   g657(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n844));
  AND2_X1   g658(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n842), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n842), .A2(new_n843), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n845), .ZN(new_n848));
  INV_X1    g662(.A(new_n728), .ZN(new_n849));
  OAI211_X1 g663(.A(G952), .B(new_n342), .C1(new_n816), .C2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n823), .A2(new_n513), .A3(new_n825), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n851), .B2(new_n633), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n818), .A2(KEYINPUT51), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n848), .B(new_n852), .C1(new_n834), .C2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n841), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n694), .A2(new_n765), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n807), .B(new_n670), .C1(new_n856), .C2(new_n759), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n507), .A2(new_n508), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n660), .A2(new_n858), .A3(new_n683), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n416), .A2(new_n418), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n733), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n649), .A2(new_n745), .A3(new_n670), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n702), .A2(new_n187), .A3(new_n751), .A4(new_n753), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n857), .A2(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n650), .B1(new_n856), .B2(new_n759), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n864), .A3(new_n774), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT114), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n755), .A2(new_n741), .A3(new_n745), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n711), .A2(new_n670), .A3(new_n807), .A4(new_n860), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n776), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n772), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n676), .A2(new_n721), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n620), .A2(new_n729), .A3(new_n737), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n634), .B1(new_n479), .B2(new_n858), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n657), .A2(new_n658), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n650), .B(new_n720), .C1(new_n856), .C2(new_n759), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n651), .A2(new_n877), .B1(new_n878), .B2(new_n663), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n874), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n715), .A2(new_n688), .A3(new_n746), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n750), .A2(new_n670), .A3(new_n681), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n698), .A2(new_n657), .A3(new_n700), .A4(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(KEYINPUT115), .A3(KEYINPUT52), .A4(new_n885), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n740), .B(new_n713), .C1(new_n606), .C2(new_n618), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n687), .B1(new_n887), .B2(new_n686), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(KEYINPUT52), .A3(new_n746), .A4(new_n885), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n715), .A2(new_n688), .A3(new_n746), .A4(new_n885), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n882), .A2(KEYINPUT53), .A3(new_n886), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  XOR2_X1   g710(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n897));
  NAND4_X1  g711(.A1(new_n725), .A2(new_n644), .A3(new_n636), .A4(new_n876), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n676), .A2(new_n726), .A3(new_n721), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n620), .A2(new_n729), .A3(new_n737), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n776), .A2(new_n869), .A3(new_n870), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n902), .A2(KEYINPUT114), .B1(new_n758), .B2(new_n771), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n903), .A3(new_n872), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n889), .A2(new_n892), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n896), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  INV_X1    g722(.A(new_n897), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n868), .A2(new_n772), .A3(new_n872), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n894), .A3(new_n886), .A4(new_n901), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n908), .A2(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n855), .B(new_n907), .C1(new_n896), .C2(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n841), .A2(new_n854), .A3(KEYINPUT120), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n812), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n418), .A2(new_n187), .ZN(new_n919));
  NOR4_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n782), .A4(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n825), .A2(new_n706), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n921), .ZN(G75));
  NAND2_X1  g736(.A1(new_n889), .A2(new_n892), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n909), .B1(new_n882), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n894), .A2(new_n886), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT53), .A4(new_n872), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(G210), .B(G902), .C1(new_n924), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n275), .A2(new_n304), .A3(new_n306), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n303), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n342), .A2(G952), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT123), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n404), .B1(new_n895), .B2(new_n906), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n933), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n928), .A2(new_n929), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(KEYINPUT122), .A3(new_n932), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n937), .B1(new_n941), .B2(new_n943), .ZN(G51));
  INV_X1    g758(.A(new_n936), .ZN(new_n945));
  NAND2_X1  g759(.A1(G469), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT57), .Z(new_n947));
  NOR3_X1   g761(.A1(new_n924), .A2(new_n927), .A3(KEYINPUT54), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n896), .B1(new_n895), .B2(new_n906), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n413), .A2(new_n414), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n939), .A2(new_n792), .A3(new_n791), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(G54));
  INV_X1    g768(.A(new_n939), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n455), .A2(new_n462), .ZN(new_n956));
  NAND2_X1  g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n945), .B1(new_n958), .B2(new_n959), .ZN(G60));
  INV_X1    g774(.A(new_n626), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n629), .B(KEYINPUT59), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n961), .B(new_n963), .C1(new_n948), .C2(new_n949), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n936), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n907), .B1(new_n913), .B2(new_n896), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n966), .B2(new_n963), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n895), .B2(new_n906), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(new_n545), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n945), .B1(new_n971), .B2(new_n668), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n971), .B2(new_n668), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n972), .B(new_n973), .C1(new_n975), .C2(KEYINPUT61), .ZN(new_n976));
  INV_X1    g790(.A(new_n970), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n668), .B(new_n977), .C1(new_n924), .C2(new_n927), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n978), .B(new_n936), .C1(new_n545), .C2(new_n971), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT61), .B1(new_n978), .B2(KEYINPUT124), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n976), .A2(new_n981), .ZN(G66));
  OAI21_X1  g796(.A(G953), .B1(new_n516), .B2(new_n299), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n901), .B2(G953), .ZN(new_n984));
  INV_X1    g798(.A(G898), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n930), .B1(new_n985), .B2(G953), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n984), .B(new_n986), .Z(G69));
  NAND2_X1  g801(.A1(new_n799), .A2(new_n809), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n843), .A2(new_n339), .A3(new_n699), .A4(new_n796), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n772), .A2(new_n883), .A3(new_n776), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n342), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n571), .A2(new_n574), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n449), .A2(new_n450), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n992), .B(new_n995), .C1(new_n680), .C2(new_n342), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n619), .A2(new_n807), .A3(new_n876), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(new_n691), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n799), .A2(new_n809), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n709), .A2(new_n883), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n709), .A2(new_n883), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT125), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT125), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n999), .A2(new_n1001), .A3(new_n1006), .A4(new_n1003), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n996), .B1(new_n1008), .B2(new_n995), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n342), .B1(G227), .B2(G900), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1010), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1012), .B(new_n996), .C1(new_n1008), .C2(new_n995), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(G72));
  NAND3_X1  g828(.A1(new_n1005), .A2(new_n901), .A3(new_n1007), .ZN(new_n1015));
  XNOR2_X1  g829(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n637), .A2(new_n404), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT127), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n695), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n611), .A2(new_n585), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n1018), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n913), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1019), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(new_n991), .B2(new_n901), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n610), .A2(new_n584), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n936), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1020), .A2(new_n1023), .A3(new_n1027), .ZN(G57));
endmodule


