//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  AND2_X1   g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n219), .B(new_n223), .C1(G107), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G238), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n218), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT68), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT69), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT70), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n213), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT15), .B(G87), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n207), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n254), .A2(new_n255), .B1(new_n207), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n253), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n263), .A2(new_n207), .A3(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n206), .A2(G20), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT74), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(new_n253), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n262), .B(new_n265), .C1(new_n269), .C2(new_n256), .ZN(new_n270));
  XOR2_X1   g0070(.A(new_n270), .B(KEYINPUT77), .Z(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G107), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n278), .B1(new_n279), .B2(new_n276), .C1(new_n281), .C2(new_n226), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT71), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(G244), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n271), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT76), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(G169), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n292), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n303), .A2(new_n271), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n264), .A2(G50), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n269), .B2(G50), .ZN(new_n307));
  INV_X1    g0107(.A(new_n253), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n258), .A2(new_n255), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n280), .A2(G223), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n276), .A2(new_n277), .ZN(new_n314));
  INV_X1    g0114(.A(G222), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(new_n256), .B2(new_n276), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n283), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n290), .A2(G226), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n285), .B(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n318), .B2(new_n320), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n317), .B(new_n326), .C1(new_n323), .C2(new_n322), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n312), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n329), .A2(KEYINPUT75), .A3(G179), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n328), .B2(new_n302), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT78), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G33), .A3(G97), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n336), .B(new_n341), .C1(new_n314), .C2(new_n235), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n283), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n286), .B1(G238), .B2(new_n290), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n343), .B2(new_n344), .ZN(new_n348));
  OAI21_X1  g0148(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT14), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(KEYINPUT79), .ZN(new_n351));
  INV_X1    g0151(.A(new_n348), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT79), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n343), .A2(new_n344), .A3(new_n353), .A4(new_n345), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n351), .A2(new_n352), .A3(G179), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n350), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT66), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT66), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n207), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n260), .A2(new_n202), .B1(new_n255), .B2(new_n256), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n253), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT11), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n225), .A2(new_n264), .A3(KEYINPUT12), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(KEYINPUT12), .B2(new_n264), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n269), .A2(KEYINPUT12), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G68), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(KEYINPUT80), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(KEYINPUT80), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n294), .B1(new_n352), .B2(new_n346), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n351), .A2(new_n352), .A3(G190), .A4(new_n354), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n358), .A2(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n305), .A2(new_n335), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n258), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n264), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n269), .B2(new_n380), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT81), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n259), .A2(G159), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n201), .B1(new_n363), .B2(G58), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(new_n207), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n274), .A2(new_n207), .A3(new_n275), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n275), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n225), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n383), .B(new_n384), .C1(new_n387), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n216), .B1(new_n225), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n396));
  AND2_X1   g0196(.A1(KEYINPUT3), .A2(G33), .ZN(new_n397));
  NOR2_X1   g0197(.A1(KEYINPUT3), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n399), .B2(new_n207), .ZN(new_n400));
  INV_X1    g0200(.A(new_n391), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n402), .A3(KEYINPUT16), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n393), .A2(new_n253), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n363), .B1(new_n400), .B2(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n383), .B1(new_n406), .B2(new_n384), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n382), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n286), .B1(G232), .B2(new_n290), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n276), .A2(G223), .A3(new_n277), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT83), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  OAI211_X1 g0213(.A(G226), .B(G1698), .C1(new_n397), .C2(new_n398), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n283), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n414), .A2(new_n413), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n417), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n410), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n294), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n297), .B(new_n410), .C1(new_n416), .C2(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  INV_X1    g0224(.A(new_n421), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT83), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n283), .A3(new_n415), .ZN(new_n428));
  AOI21_X1  g0228(.A(G200), .B1(new_n428), .B2(new_n410), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n382), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n393), .A2(new_n253), .A3(new_n403), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n407), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n424), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT82), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT82), .B(new_n431), .C1(new_n432), .C2(new_n407), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n419), .A2(new_n330), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n428), .A2(new_n302), .A3(new_n410), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT18), .A4(new_n441), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n435), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n325), .A2(G200), .A3(new_n327), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT9), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n312), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n297), .B1(new_n325), .B2(new_n327), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT10), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n328), .A2(G190), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT10), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n447), .A4(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n379), .A2(new_n446), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G283), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n273), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n280), .B2(G250), .ZN(new_n460));
  OAI211_X1 g0260(.A(G244), .B(new_n277), .C1(new_n397), .C2(new_n398), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT86), .A2(KEYINPUT4), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT86), .A2(KEYINPUT4), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n461), .B2(new_n462), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n283), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n288), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(new_n213), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G41), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n206), .A2(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n472), .A2(G257), .B1(G274), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n467), .A2(new_n297), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n467), .A2(new_n478), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(G200), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n279), .A2(KEYINPUT6), .A3(G97), .ZN(new_n482));
  AND2_X1   g0282(.A1(G97), .A2(G107), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n482), .B1(new_n485), .B2(KEYINPUT6), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n487));
  OAI21_X1  g0287(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n308), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n264), .A2(new_n221), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT85), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n268), .B1(G1), .B2(new_n273), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n481), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n207), .B(G87), .C1(new_n397), .C2(new_n398), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n276), .A2(new_n501), .A3(new_n207), .A4(G87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT91), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n207), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n279), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n504), .B1(new_n503), .B2(new_n510), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n498), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n503), .A2(new_n510), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT24), .A3(new_n511), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n517), .A3(new_n253), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n263), .A2(G1), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(G20), .A3(new_n279), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT25), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n495), .B2(G107), .ZN(new_n522));
  OAI211_X1 g0322(.A(G250), .B(new_n277), .C1(new_n397), .C2(new_n398), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(G1698), .C1(new_n397), .C2(new_n398), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G294), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n283), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n472), .A2(KEYINPUT92), .A3(G264), .ZN(new_n528));
  AND2_X1   g0328(.A1(KEYINPUT5), .A2(G41), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n469), .B1(new_n529), .B2(new_n474), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n470), .A2(new_n471), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(G264), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT92), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n477), .A2(G274), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n527), .A2(new_n528), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n294), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G190), .B2(new_n536), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n518), .A2(new_n522), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n467), .A2(G179), .A3(new_n478), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n480), .B2(new_n330), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n543), .B(new_n308), .C1(new_n487), .C2(new_n488), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n496), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n473), .A2(G250), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n469), .A2(G274), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n283), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G238), .B(new_n277), .C1(new_n397), .C2(new_n398), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(G1698), .C1(new_n397), .C2(new_n398), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n505), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(new_n283), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n294), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n338), .B2(new_n340), .ZN(new_n556));
  INV_X1    g0356(.A(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n221), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n556), .A2(G20), .B1(G107), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(G20), .B1(new_n274), .B2(new_n275), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(G68), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n308), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n254), .ZN(new_n564));
  INV_X1    g0364(.A(new_n264), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n494), .A2(new_n557), .ZN(new_n567));
  NOR4_X1   g0367(.A1(new_n554), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n552), .A2(new_n283), .ZN(new_n570));
  INV_X1    g0370(.A(new_n549), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n297), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n553), .A2(KEYINPUT87), .A3(G190), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n563), .A2(new_n566), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n254), .B2(new_n494), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n553), .A2(G179), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n330), .B2(new_n553), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n568), .A2(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n497), .A2(new_n539), .A3(new_n546), .A4(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT21), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n565), .A2(G116), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n495), .B2(G116), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(G20), .B1(new_n273), .B2(G97), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n273), .B2(new_n458), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  INV_X1    g0389(.A(G116), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G20), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n253), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n253), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT90), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT20), .B(new_n588), .C1(new_n592), .C2(new_n593), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT89), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n586), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n472), .A2(G270), .B1(G274), .B2(new_n477), .ZN(new_n605));
  OAI211_X1 g0405(.A(G264), .B(G1698), .C1(new_n397), .C2(new_n398), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n277), .C1(new_n397), .C2(new_n398), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n274), .A2(G303), .A3(new_n275), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n283), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n330), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n583), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n599), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n597), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(KEYINPUT21), .A3(G169), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n605), .A2(new_n610), .A3(G179), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n619), .A2(new_n585), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n611), .A2(new_n294), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G190), .B2(new_n611), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n604), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n615), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n518), .A2(new_n522), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n536), .A2(G169), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n302), .B2(new_n536), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n582), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n457), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT93), .ZN(G372));
  NAND2_X1  g0435(.A1(new_n619), .A2(new_n585), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n613), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n622), .B1(new_n637), .B2(new_n583), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n631), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n582), .B1(new_n577), .B2(new_n579), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n568), .A2(new_n575), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n577), .A2(new_n579), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n545), .A2(new_n641), .A3(new_n541), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n580), .A2(new_n545), .A3(new_n541), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n457), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n335), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n441), .A2(new_n433), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT18), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n441), .A2(new_n433), .A3(new_n443), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n358), .A2(new_n374), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n304), .A2(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n303), .A2(new_n271), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT94), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n376), .A2(new_n377), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n655), .B1(new_n664), .B2(new_n435), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT95), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n452), .A2(new_n666), .A3(new_n455), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n452), .B2(new_n455), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n650), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n649), .A2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n519), .A2(new_n207), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n638), .A2(new_n636), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n677), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n604), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n627), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT96), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT97), .B(G330), .Z(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n628), .A2(new_n630), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n628), .A2(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n539), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n631), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n682), .A2(new_n684), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n686), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n615), .A2(new_n623), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n679), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n686), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n690), .A2(new_n696), .ZN(G399));
  NAND2_X1  g0497(.A1(new_n210), .A2(new_n287), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n558), .A2(G107), .A3(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n218), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n648), .A2(new_n679), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT102), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n644), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n647), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT102), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n677), .B1(new_n710), .B2(new_n640), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n528), .A2(new_n534), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(KEYINPUT98), .A3(new_n527), .A4(new_n553), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT98), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n572), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n621), .A2(KEYINPUT99), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT99), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n605), .A2(new_n610), .A3(new_n721), .A4(G179), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n719), .A2(KEYINPUT30), .A3(new_n480), .A4(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n612), .A2(G179), .A3(new_n553), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n467), .A2(new_n478), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n536), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n715), .B2(new_n718), .ZN(new_n730));
  AOI211_X1 g0530(.A(KEYINPUT101), .B(KEYINPUT30), .C1(new_n730), .C2(new_n723), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT101), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT98), .B1(new_n733), .B2(new_n553), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n717), .A2(new_n572), .A3(new_n716), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n723), .B(new_n480), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n728), .B(new_n729), .C1(new_n731), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n677), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n631), .A2(new_n615), .A3(new_n623), .A4(new_n626), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT31), .B1(new_n741), .B2(new_n581), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n679), .A2(new_n729), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n724), .A2(new_n727), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT30), .B1(new_n730), .B2(new_n723), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT100), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n683), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n713), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n702), .B1(new_n753), .B2(G1), .ZN(G364));
  OR2_X1    g0554(.A1(new_n682), .A2(new_n684), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n682), .A2(new_n684), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n263), .A2(G20), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G45), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n698), .A2(G1), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n213), .B1(G20), .B2(new_n330), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n302), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n207), .B1(new_n766), .B2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n764), .A2(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(new_n297), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n302), .A2(new_n294), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT103), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n772), .A2(KEYINPUT103), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n769), .B1(new_n777), .B2(G326), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT104), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n770), .A2(new_n763), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n276), .B1(new_n781), .B2(G322), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n294), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n770), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n762), .A2(new_n766), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G303), .A2(new_n785), .B1(new_n787), .B2(G329), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n771), .A2(new_n762), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n762), .A2(new_n783), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n790), .A2(new_n791), .B1(new_n793), .B2(G283), .ZN(new_n794));
  AND4_X1   g0594(.A1(new_n779), .A2(new_n782), .A3(new_n788), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n786), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n202), .B2(new_n776), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G68), .A2(new_n790), .B1(new_n793), .B2(G107), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n800), .B1(new_n394), .B2(new_n780), .C1(new_n557), .C2(new_n784), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n276), .B1(new_n767), .B2(new_n221), .C1(new_n256), .C2(new_n764), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n761), .B1(new_n795), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n761), .ZN(new_n808));
  INV_X1    g0608(.A(new_n210), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n276), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n247), .A2(new_n288), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n218), .A2(new_n288), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n210), .A2(new_n276), .ZN(new_n815));
  INV_X1    g0615(.A(G355), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n816), .B1(G116), .B2(new_n210), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n808), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n759), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n804), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n681), .B2(new_n807), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n760), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NAND4_X1  g0623(.A1(new_n658), .A2(new_n271), .A3(new_n661), .A4(new_n677), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n271), .A2(new_n677), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n659), .B(new_n825), .C1(new_n296), .C2(new_n299), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n703), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n751), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n819), .B1(new_n828), .B2(new_n751), .ZN(new_n831));
  INV_X1    g0631(.A(new_n827), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n805), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n789), .A2(new_n458), .B1(new_n764), .B2(new_n590), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n777), .B2(G303), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT105), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n399), .B1(new_n780), .B2(new_n768), .ZN(new_n837));
  INV_X1    g0637(.A(new_n767), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(G97), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G107), .A2(new_n785), .B1(new_n793), .B2(G87), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n839), .B(new_n840), .C1(new_n765), .C2(new_n786), .ZN(new_n841));
  INV_X1    g0641(.A(new_n764), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G150), .A2(new_n790), .B1(new_n842), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G143), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n844), .B2(new_n780), .C1(new_n776), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(KEYINPUT34), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n276), .B1(new_n784), .B2(new_n202), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n792), .A2(new_n359), .B1(new_n786), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(G58), .C2(new_n838), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n836), .A2(new_n841), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(new_n761), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n761), .A2(new_n805), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n759), .B(new_n856), .C1(new_n256), .C2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n830), .A2(new_n831), .B1(new_n833), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  OAI21_X1  g0660(.A(G77), .B1(new_n225), .B2(new_n394), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n218), .A2(new_n861), .B1(G50), .B2(new_n359), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(G1), .A3(new_n263), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT106), .Z(new_n864));
  OAI211_X1 g0664(.A(G116), .B(new_n214), .C1(new_n486), .C2(KEYINPUT35), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(KEYINPUT35), .B2(new_n486), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT36), .Z(new_n867));
  OAI21_X1  g0667(.A(new_n728), .B1(new_n731), .B2(new_n738), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n740), .A2(new_n742), .B1(new_n868), .B2(new_n745), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n374), .A2(new_n677), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n657), .A2(new_n677), .B1(new_n378), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n869), .A2(new_n832), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n675), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n437), .A2(new_n438), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT37), .B1(new_n409), .B2(new_n422), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n442), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n439), .A2(new_n440), .ZN(new_n877));
  INV_X1    g0677(.A(new_n402), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n384), .B1(new_n878), .B2(new_n387), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n403), .A3(new_n253), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n877), .A2(new_n675), .B1(new_n880), .B2(new_n431), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n430), .A2(new_n433), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n431), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n873), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n446), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n884), .C1(new_n446), .C2(new_n886), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n872), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n437), .A2(new_n438), .A3(new_n873), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n409), .A2(new_n422), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n651), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n876), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n654), .B2(new_n435), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n888), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n893), .B1(new_n901), .B2(new_n890), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n892), .A2(new_n893), .B1(new_n872), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n868), .A2(new_n745), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n743), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n457), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n903), .B(new_n906), .Z(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(new_n683), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n692), .A2(new_n685), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n642), .B1(new_n909), .B2(new_n581), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n644), .A2(new_n647), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n827), .B(new_n679), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n659), .A2(new_n677), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n871), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n891), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n654), .A2(new_n675), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT107), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n898), .B2(new_n899), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n889), .B(new_n890), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT39), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n901), .A2(new_n890), .ZN(new_n923));
  NOR2_X1   g0723(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n656), .A2(new_n677), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n705), .A2(new_n712), .A3(new_n457), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n670), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n908), .A2(new_n931), .B1(new_n206), .B2(new_n757), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n908), .A2(new_n931), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n864), .B(new_n867), .C1(new_n932), .C2(new_n933), .ZN(G367));
  INV_X1    g0734(.A(new_n761), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n777), .A2(G143), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n789), .A2(new_n796), .B1(new_n792), .B2(new_n256), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n399), .B(new_n937), .C1(G137), .C2(new_n787), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n838), .A2(G68), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n784), .A2(new_n394), .B1(new_n764), .B2(new_n202), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G150), .B2(new_n781), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n936), .A2(new_n938), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n777), .A2(G311), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n792), .A2(new_n221), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n784), .A2(new_n590), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n276), .B(new_n944), .C1(KEYINPUT46), .C2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(KEYINPUT46), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G107), .B2(new_n838), .ZN(new_n948));
  INV_X1    g0748(.A(G303), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n780), .A2(new_n949), .B1(new_n764), .B2(new_n458), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n789), .A2(new_n768), .B1(new_n786), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n943), .A2(new_n946), .A3(new_n948), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n942), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT109), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT47), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n935), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n242), .A2(new_n810), .ZN(new_n960));
  INV_X1    g0760(.A(new_n808), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n809), .B2(new_n564), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n759), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n807), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n495), .A2(G87), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n679), .B1(new_n576), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n580), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n642), .B2(new_n966), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n959), .B(new_n963), .C1(new_n964), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n758), .A2(G1), .ZN(new_n970));
  INV_X1    g0770(.A(new_n690), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n545), .A2(new_n677), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n497), .A2(new_n546), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n541), .A2(new_n545), .A3(new_n677), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n696), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n696), .A2(KEYINPUT44), .A3(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT44), .B1(new_n696), .B2(new_n975), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n971), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n976), .B(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n983), .A2(new_n690), .A3(new_n979), .A4(new_n978), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n682), .A2(KEYINPUT108), .A3(new_n684), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n691), .B(new_n693), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT108), .B1(new_n682), .B2(new_n684), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n753), .B1(new_n985), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n698), .B(KEYINPUT41), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n970), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n694), .A2(new_n975), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n546), .B1(new_n973), .B2(new_n631), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n679), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n690), .B1(new_n974), .B2(new_n973), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n969), .B1(new_n996), .B2(new_n1009), .ZN(G387));
  NAND2_X1  g0810(.A1(new_n993), .A2(new_n752), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n992), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n990), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n753), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n698), .B(KEYINPUT111), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n815), .A2(new_n699), .B1(G107), .B2(new_n210), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n238), .A2(G45), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n699), .ZN(new_n1019));
  AOI211_X1 g0819(.A(G45), .B(new_n1019), .C1(G68), .C2(G77), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n258), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n811), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1017), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n819), .B1(new_n1024), .B2(new_n961), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G317), .A2(new_n781), .B1(new_n842), .B2(G303), .ZN(new_n1026));
  INV_X1    g0826(.A(G322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n765), .B2(new_n789), .C1(new_n776), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n785), .A2(G294), .B1(new_n838), .B2(G283), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n399), .B1(new_n792), .B2(new_n590), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G326), .B2(new_n787), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(G150), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n789), .A2(new_n258), .B1(new_n786), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G77), .B2(new_n785), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n780), .A2(new_n202), .B1(new_n764), .B2(new_n359), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n767), .A2(new_n254), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1043), .A2(new_n944), .A3(new_n1044), .A4(new_n399), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT110), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n777), .B2(G159), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n776), .A2(KEYINPUT110), .A3(new_n796), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1042), .B(new_n1045), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n935), .B1(new_n1039), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1025), .B(new_n1050), .C1(new_n691), .C2(new_n807), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1013), .B2(new_n970), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1016), .A2(new_n1052), .ZN(G393));
  NAND2_X1  g0853(.A1(new_n810), .A2(new_n250), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n808), .C1(new_n221), .C2(new_n210), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT112), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n819), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n776), .A2(new_n1040), .B1(new_n796), .B2(new_n780), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n276), .B1(new_n767), .B2(new_n256), .C1(new_n557), .C2(new_n792), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n789), .A2(new_n202), .B1(new_n764), .B2(new_n258), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n784), .A2(new_n225), .B1(new_n786), .B2(new_n844), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n776), .A2(new_n951), .B1(new_n765), .B2(new_n780), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n399), .B1(new_n767), .B2(new_n590), .C1(new_n279), .C2(new_n792), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n784), .A2(new_n458), .B1(new_n786), .B2(new_n1027), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n789), .A2(new_n949), .B1(new_n764), .B2(new_n768), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1061), .A2(new_n1065), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT113), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n935), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1059), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n964), .B2(new_n975), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n970), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n985), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1015), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n981), .A2(new_n984), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n752), .B1(new_n990), .B2(new_n1012), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1014), .A2(new_n985), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1079), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  AOI21_X1  g0886(.A(new_n759), .B1(new_n258), .B2(new_n857), .ZN(new_n1087));
  INV_X1    g0887(.A(G128), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n776), .A2(new_n1088), .B1(new_n850), .B2(new_n780), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT115), .Z(new_n1090));
  NAND2_X1  g0890(.A1(new_n785), .A2(G150), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT53), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G50), .A2(new_n793), .B1(new_n787), .B2(G125), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n764), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n276), .B1(new_n767), .B2(new_n796), .C1(new_n845), .C2(new_n789), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n399), .B1(new_n784), .B2(new_n557), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n789), .A2(new_n279), .B1(new_n792), .B2(new_n359), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G77), .C2(new_n838), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G116), .A2(new_n781), .B1(new_n787), .B2(G294), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n221), .B2(new_n764), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G283), .B2(new_n777), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1090), .A2(new_n1097), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1087), .B1(new_n935), .B2(new_n1104), .C1(new_n926), .C2(new_n806), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(KEYINPUT39), .A2(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n927), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n912), .A2(new_n914), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n871), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n923), .A2(new_n927), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n913), .B1(new_n711), .B2(new_n827), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n871), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n684), .B(new_n827), .C1(new_n744), .C2(new_n749), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(new_n871), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1110), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1112), .A2(new_n871), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1106), .A2(new_n1109), .B1(new_n1117), .B2(new_n1111), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n869), .A2(new_n832), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n871), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(G330), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1116), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1105), .B1(new_n1122), .B2(new_n1078), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1110), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n457), .A2(G330), .A3(new_n905), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n929), .A2(new_n670), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT114), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n929), .A2(KEYINPUT114), .A3(new_n670), .A4(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1112), .B1(new_n871), .B2(new_n1114), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1120), .B1(new_n1119), .B2(G330), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1114), .A2(new_n871), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1108), .B1(new_n1136), .B2(new_n1121), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1080), .B1(new_n1126), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1122), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1123), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(G378));
  INV_X1    g0944(.A(new_n1132), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1122), .B2(new_n1138), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n916), .B(new_n917), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n889), .A2(new_n890), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n905), .A2(new_n827), .A3(new_n1120), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n893), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n873), .B1(new_n307), .B2(new_n311), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT55), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n669), .B2(new_n335), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n456), .A2(KEYINPUT95), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n452), .A2(new_n455), .A3(new_n666), .ZN(new_n1157));
  AND4_X1   g0957(.A1(new_n335), .A2(new_n1156), .A3(new_n1157), .A4(new_n1154), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1153), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n669), .A2(new_n335), .A3(new_n1154), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1156), .A2(new_n335), .A3(new_n1157), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1154), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1160), .A2(new_n1163), .A3(new_n1152), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n902), .A2(new_n872), .ZN(new_n1166));
  AND4_X1   g0966(.A1(G330), .A2(new_n1150), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n903), .B2(G330), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1147), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1150), .A2(G330), .A3(new_n1166), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1165), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n903), .A2(G330), .A3(new_n1165), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n928), .A3(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1146), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1176), .B1(new_n1146), .B2(new_n1175), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1015), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1169), .A2(new_n970), .A3(new_n1174), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n759), .B1(new_n202), .B2(new_n857), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n764), .A2(new_n254), .B1(new_n786), .B2(new_n458), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G107), .B2(new_n781), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n256), .A2(new_n784), .B1(new_n789), .B2(new_n221), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n792), .A2(new_n394), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n399), .A2(new_n287), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n939), .B1(new_n776), .B2(new_n590), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT117), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1183), .B(new_n1187), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n780), .A2(new_n1088), .B1(new_n764), .B2(new_n845), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n850), .A2(new_n789), .B1(new_n784), .B2(new_n1094), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G150), .C2(new_n838), .ZN(new_n1197));
  INV_X1    g0997(.A(G125), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n776), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n273), .B(new_n287), .C1(new_n792), .C2(new_n796), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G124), .B2(new_n787), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1186), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT116), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1194), .A2(new_n1204), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1181), .B1(new_n935), .B2(new_n1208), .C1(new_n1171), .C2(new_n806), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1180), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1179), .A2(new_n1211), .ZN(G375));
  AOI21_X1  g1012(.A(new_n759), .B1(new_n359), .B2(new_n857), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n590), .A2(new_n789), .B1(new_n780), .B2(new_n458), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n399), .B1(new_n792), .B2(new_n256), .ZN(new_n1215));
  OR3_X1    g1015(.A1(new_n1214), .A2(new_n1044), .A3(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G97), .A2(new_n785), .B1(new_n787), .B2(G303), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n279), .B2(new_n764), .C1(new_n776), .C2(new_n768), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G159), .A2(new_n785), .B1(new_n787), .B2(G128), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n1040), .B2(new_n764), .C1(new_n776), .C2(new_n850), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n845), .A2(new_n780), .B1(new_n789), .B2(new_n1094), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n767), .A2(new_n202), .ZN(new_n1222));
  OR4_X1    g1022(.A1(new_n399), .A2(new_n1221), .A3(new_n1185), .A4(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1216), .A2(new_n1218), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT119), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n761), .B1(new_n1224), .B2(KEYINPUT119), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1213), .B1(new_n1225), .B2(new_n1226), .C1(new_n1120), .C2(new_n806), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1138), .B2(new_n1078), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1141), .A2(new_n995), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1138), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1145), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1229), .B1(new_n1230), .B2(new_n1232), .ZN(G381));
  NAND3_X1  g1033(.A1(new_n1016), .A2(new_n822), .A3(new_n1052), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT120), .B1(new_n1235), .B2(new_n859), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1085), .B(new_n969), .C1(new_n996), .C2(new_n1009), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT120), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1234), .A2(new_n1238), .A3(G384), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .A4(G381), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT121), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1179), .A2(new_n1143), .A3(new_n1211), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1241), .A2(new_n1242), .ZN(G407));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G343), .C2(new_n1242), .ZN(G409));
  INV_X1    g1044(.A(G213), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(G343), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1210), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1146), .A2(new_n1175), .A3(new_n995), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1180), .A2(KEYINPUT122), .A3(new_n1209), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1143), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1251), .B2(new_n1143), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1179), .A2(G378), .A3(new_n1211), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1246), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1232), .A2(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1145), .A2(new_n1231), .A3(KEYINPUT60), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1015), .B(new_n1141), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(G384), .A3(new_n1229), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G384), .B1(new_n1261), .B2(new_n1229), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G2897), .B(new_n1246), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(G2897), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1262), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT63), .B1(new_n1257), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1251), .A2(new_n1143), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT123), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1251), .A2(new_n1143), .A3(new_n1252), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1256), .A3(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1246), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1257), .A2(KEYINPUT63), .A3(new_n1275), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(G390), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1237), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT126), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n822), .B1(new_n1016), .B2(new_n1052), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT124), .B1(new_n1235), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1284), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1234), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1280), .A2(new_n1290), .A3(new_n1237), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1283), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1289), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT126), .A3(new_n1282), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(KEYINPUT61), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1278), .A2(new_n1279), .A3(new_n1296), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1277), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1257), .B2(new_n1269), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1277), .B2(KEYINPUT127), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1295), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1297), .B1(new_n1302), .B2(new_n1303), .ZN(G405));
  AND3_X1   g1104(.A1(new_n1292), .A2(new_n1294), .A3(new_n1275), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1275), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(G375), .B(new_n1143), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1307), .B(new_n1308), .ZN(G402));
endmodule


