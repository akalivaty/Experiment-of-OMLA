

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782;

  INV_X2 U381 ( .A(G953), .ZN(n768) );
  AND2_X1 U382 ( .A1(n431), .A2(n568), .ZN(n424) );
  INV_X1 U383 ( .A(n673), .ZN(n767) );
  BUF_X1 U384 ( .A(n747), .Z(n360) );
  AND2_X4 U385 ( .A1(n442), .A2(n443), .ZN(n747) );
  XNOR2_X2 U386 ( .A(n412), .B(n484), .ZN(n507) );
  XNOR2_X2 U387 ( .A(G119), .B(KEYINPUT70), .ZN(n392) );
  XNOR2_X2 U388 ( .A(n489), .B(G469), .ZN(n597) );
  NOR2_X1 U389 ( .A1(n573), .A2(n556), .ZN(n557) );
  AND2_X1 U390 ( .A1(n564), .A2(n563), .ZN(n653) );
  XNOR2_X1 U391 ( .A(n619), .B(n618), .ZN(n388) );
  AND2_X1 U392 ( .A1(n385), .A2(n384), .ZN(n579) );
  NAND2_X1 U393 ( .A1(n380), .A2(n387), .ZN(n720) );
  AND2_X1 U394 ( .A1(n393), .A2(n705), .ZN(n617) );
  AND2_X1 U395 ( .A1(n381), .A2(n457), .ZN(n380) );
  XNOR2_X1 U396 ( .A(n693), .B(n458), .ZN(n603) );
  XNOR2_X1 U397 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U398 ( .A(n437), .B(n506), .ZN(n685) );
  NAND2_X1 U399 ( .A1(n378), .A2(n410), .ZN(n409) );
  XNOR2_X1 U400 ( .A(n740), .B(n479), .ZN(n741) );
  XNOR2_X1 U401 ( .A(n539), .B(n430), .ZN(n740) );
  XNOR2_X1 U402 ( .A(G143), .B(G128), .ZN(n517) );
  XNOR2_X1 U403 ( .A(n392), .B(n391), .ZN(n390) );
  XNOR2_X1 U404 ( .A(n390), .B(n389), .ZN(n377) );
  BUF_X1 U405 ( .A(n757), .Z(n361) );
  XNOR2_X1 U406 ( .A(n377), .B(n516), .ZN(n757) );
  BUF_X1 U407 ( .A(n640), .Z(n441) );
  BUF_X1 U408 ( .A(n642), .Z(n752) );
  XOR2_X1 U409 ( .A(KEYINPUT4), .B(G101), .Z(n510) );
  XNOR2_X1 U410 ( .A(n480), .B(G116), .ZN(n389) );
  INV_X1 U411 ( .A(G113), .ZN(n480) );
  XNOR2_X1 U412 ( .A(G902), .B(KEYINPUT15), .ZN(n518) );
  NAND2_X1 U413 ( .A1(n402), .A2(n401), .ZN(n400) );
  INV_X1 U414 ( .A(n409), .ZN(n402) );
  NOR2_X1 U415 ( .A1(n362), .A2(n365), .ZN(n401) );
  AND2_X1 U416 ( .A1(n405), .A2(n371), .ZN(n403) );
  NAND2_X1 U417 ( .A1(n409), .A2(n406), .ZN(n405) );
  OR2_X1 U418 ( .A1(n365), .A2(n704), .ZN(n404) );
  XNOR2_X1 U419 ( .A(n558), .B(n386), .ZN(n385) );
  INV_X1 U420 ( .A(KEYINPUT22), .ZN(n386) );
  NOR2_X1 U421 ( .A1(n620), .A2(n686), .ZN(n460) );
  OR2_X2 U422 ( .A1(n362), .A2(n409), .ZN(n693) );
  NAND2_X1 U423 ( .A1(n566), .A2(n473), .ZN(n470) );
  NOR2_X1 U424 ( .A1(n465), .A2(n464), .ZN(n463) );
  NAND2_X1 U425 ( .A1(n633), .A2(n363), .ZN(n396) );
  INV_X1 U426 ( .A(KEYINPUT48), .ZN(n395) );
  NOR2_X1 U427 ( .A1(n581), .A2(n582), .ZN(n583) );
  NAND2_X1 U428 ( .A1(n399), .A2(n406), .ZN(n398) );
  INV_X1 U429 ( .A(n407), .ZN(n399) );
  XNOR2_X1 U430 ( .A(n517), .B(G134), .ZN(n547) );
  XNOR2_X1 U431 ( .A(n547), .B(n451), .ZN(n764) );
  XNOR2_X1 U432 ( .A(n531), .B(n452), .ZN(n451) );
  XNOR2_X1 U433 ( .A(n453), .B(G137), .ZN(n452) );
  INV_X1 U434 ( .A(KEYINPUT68), .ZN(n453) );
  XNOR2_X1 U435 ( .A(n517), .B(n514), .ZN(n419) );
  XOR2_X1 U436 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n509) );
  XNOR2_X1 U437 ( .A(n759), .B(n474), .ZN(n512) );
  INV_X1 U438 ( .A(KEYINPUT71), .ZN(n474) );
  NOR2_X1 U439 ( .A1(n689), .A2(KEYINPUT33), .ZN(n455) );
  XNOR2_X1 U440 ( .A(n520), .B(n519), .ZN(n640) );
  NAND2_X1 U441 ( .A1(n411), .A2(G902), .ZN(n410) );
  XNOR2_X1 U442 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U443 ( .A(KEYINPUT25), .ZN(n504) );
  XNOR2_X1 U444 ( .A(G122), .B(KEYINPUT16), .ZN(n516) );
  XNOR2_X1 U445 ( .A(n476), .B(n475), .ZN(n759) );
  XNOR2_X1 U446 ( .A(G110), .B(KEYINPUT76), .ZN(n475) );
  XNOR2_X1 U447 ( .A(n477), .B(G104), .ZN(n476) );
  INV_X1 U448 ( .A(G107), .ZN(n477) );
  XNOR2_X1 U449 ( .A(n454), .B(G131), .ZN(n531) );
  INV_X1 U450 ( .A(KEYINPUT67), .ZN(n454) );
  XNOR2_X1 U451 ( .A(n494), .B(n513), .ZN(n766) );
  XNOR2_X1 U452 ( .A(n429), .B(n485), .ZN(n494) );
  XNOR2_X1 U453 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n429) );
  NOR2_X1 U454 ( .A1(G953), .A2(G237), .ZN(n481) );
  XNOR2_X1 U455 ( .A(G143), .B(G122), .ZN(n532) );
  AND2_X1 U456 ( .A1(n752), .A2(n427), .ZN(n672) );
  NOR2_X1 U457 ( .A1(n673), .A2(n428), .ZN(n427) );
  INV_X1 U458 ( .A(KEYINPUT2), .ZN(n428) );
  INV_X1 U459 ( .A(KEYINPUT84), .ZN(n439) );
  XNOR2_X1 U460 ( .A(n543), .B(n542), .ZN(n573) );
  XNOR2_X1 U461 ( .A(n541), .B(G475), .ZN(n542) );
  INV_X1 U462 ( .A(KEYINPUT87), .ZN(n423) );
  INV_X1 U463 ( .A(n685), .ZN(n440) );
  INV_X1 U464 ( .A(n603), .ZN(n384) );
  NOR2_X1 U465 ( .A1(n566), .A2(n473), .ZN(n472) );
  INV_X1 U466 ( .A(n563), .ZN(n465) );
  INV_X1 U467 ( .A(n472), .ZN(n464) );
  XNOR2_X1 U468 ( .A(n446), .B(n623), .ZN(n445) );
  AND2_X1 U469 ( .A1(n704), .A2(n365), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n508), .A2(n408), .ZN(n407) );
  INV_X1 U471 ( .A(G902), .ZN(n408) );
  XOR2_X1 U472 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n535) );
  XNOR2_X1 U473 ( .A(G113), .B(G104), .ZN(n534) );
  XOR2_X1 U474 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n533) );
  XNOR2_X1 U475 ( .A(n396), .B(n395), .ZN(n394) );
  INV_X1 U476 ( .A(n668), .ZN(n636) );
  XNOR2_X1 U477 ( .A(n421), .B(n584), .ZN(n642) );
  XOR2_X1 U478 ( .A(KEYINPUT85), .B(KEYINPUT45), .Z(n584) );
  NAND2_X1 U479 ( .A1(G234), .A2(G237), .ZN(n523) );
  XNOR2_X1 U480 ( .A(n459), .B(KEYINPUT104), .ZN(n458) );
  XNOR2_X1 U481 ( .A(n413), .B(n764), .ZN(n412) );
  XNOR2_X1 U482 ( .A(G119), .B(G137), .ZN(n495) );
  XNOR2_X1 U483 ( .A(G116), .B(G107), .ZN(n544) );
  XOR2_X1 U484 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n545) );
  XNOR2_X1 U485 ( .A(n764), .B(n366), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n417), .B(n416), .ZN(n728) );
  XNOR2_X1 U487 ( .A(n515), .B(n512), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n757), .B(n418), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n448), .B(n447), .ZN(n721) );
  INV_X1 U490 ( .A(KEYINPUT41), .ZN(n447) );
  NOR2_X1 U491 ( .A1(n701), .A2(n620), .ZN(n448) );
  AND2_X1 U492 ( .A1(n435), .A2(n614), .ZN(n393) );
  INV_X1 U493 ( .A(n615), .ZN(n436) );
  NAND2_X1 U494 ( .A1(n403), .A2(n400), .ZN(n616) );
  XNOR2_X1 U495 ( .A(n522), .B(KEYINPUT19), .ZN(n598) );
  NOR2_X1 U496 ( .A1(n640), .A2(n602), .ZN(n522) );
  AND2_X1 U497 ( .A1(n385), .A2(n690), .ZN(n561) );
  XNOR2_X1 U498 ( .A(n507), .B(KEYINPUT62), .ZN(n644) );
  XNOR2_X1 U499 ( .A(n538), .B(n370), .ZN(n430) );
  NAND2_X1 U500 ( .A1(n444), .A2(n376), .ZN(n442) );
  NOR2_X1 U501 ( .A1(G952), .A2(n768), .ZN(n751) );
  XNOR2_X1 U502 ( .A(KEYINPUT42), .B(n622), .ZN(n782) );
  NAND2_X1 U503 ( .A1(n721), .A2(n621), .ZN(n622) );
  INV_X1 U504 ( .A(n698), .ZN(n415) );
  XNOR2_X1 U505 ( .A(n580), .B(KEYINPUT106), .ZN(n777) );
  NAND2_X1 U506 ( .A1(n426), .A2(n368), .ZN(n580) );
  NOR2_X1 U507 ( .A1(n507), .A2(n407), .ZN(n362) );
  AND2_X1 U508 ( .A1(n445), .A2(n373), .ZN(n363) );
  AND2_X1 U509 ( .A1(n603), .A2(n455), .ZN(n364) );
  XOR2_X1 U510 ( .A(n613), .B(KEYINPUT111), .Z(n365) );
  XOR2_X1 U511 ( .A(G146), .B(n510), .Z(n366) );
  XNOR2_X1 U512 ( .A(n554), .B(KEYINPUT109), .ZN(n367) );
  AND2_X1 U513 ( .A1(n690), .A2(n440), .ZN(n368) );
  AND2_X1 U514 ( .A1(n636), .A2(n669), .ZN(n369) );
  AND2_X1 U515 ( .A1(G214), .A2(n540), .ZN(n370) );
  NAND2_X1 U516 ( .A1(n394), .A2(n369), .ZN(n673) );
  AND2_X1 U517 ( .A1(n397), .A2(n404), .ZN(n371) );
  AND2_X1 U518 ( .A1(n471), .A2(n470), .ZN(n372) );
  INV_X1 U519 ( .A(G140), .ZN(n485) );
  AND2_X1 U520 ( .A1(n611), .A2(n667), .ZN(n373) );
  XNOR2_X1 U521 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n374) );
  XNOR2_X1 U522 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n375) );
  NAND2_X1 U523 ( .A1(n585), .A2(KEYINPUT2), .ZN(n376) );
  INV_X1 U524 ( .A(KEYINPUT65), .ZN(n473) );
  XNOR2_X1 U525 ( .A(n377), .B(n366), .ZN(n413) );
  NAND2_X1 U526 ( .A1(n507), .A2(n411), .ZN(n378) );
  XNOR2_X1 U527 ( .A(n379), .B(n374), .ZN(n450) );
  NAND2_X1 U528 ( .A1(n383), .A2(n720), .ZN(n379) );
  NAND2_X1 U529 ( .A1(n364), .A2(n382), .ZN(n381) );
  INV_X1 U530 ( .A(n690), .ZN(n382) );
  INV_X1 U531 ( .A(n571), .ZN(n383) );
  XNOR2_X1 U532 ( .A(n461), .B(KEYINPUT93), .ZN(n571) );
  AND2_X1 U533 ( .A1(n469), .A2(n372), .ZN(n468) );
  NAND2_X1 U534 ( .A1(n414), .A2(KEYINPUT33), .ZN(n387) );
  NAND2_X1 U535 ( .A1(n579), .A2(n559), .ZN(n422) );
  XNOR2_X2 U536 ( .A(n597), .B(KEYINPUT1), .ZN(n690) );
  XNOR2_X1 U537 ( .A(n488), .B(n425), .ZN(n734) );
  NAND2_X1 U538 ( .A1(n388), .A2(n782), .ZN(n446) );
  XNOR2_X1 U539 ( .A(n388), .B(G131), .ZN(G33) );
  XNOR2_X2 U540 ( .A(KEYINPUT3), .B(KEYINPUT69), .ZN(n391) );
  NAND2_X1 U541 ( .A1(n393), .A2(n367), .ZN(n624) );
  OR2_X1 U542 ( .A1(n507), .A2(n398), .ZN(n397) );
  INV_X1 U543 ( .A(n508), .ZN(n411) );
  NAND2_X1 U544 ( .A1(n456), .A2(n603), .ZN(n414) );
  AND2_X1 U545 ( .A1(n461), .A2(n415), .ZN(n570) );
  XNOR2_X2 U546 ( .A(n462), .B(KEYINPUT0), .ZN(n461) );
  NAND2_X1 U547 ( .A1(n728), .A2(n518), .ZN(n520) );
  XNOR2_X1 U548 ( .A(n511), .B(n419), .ZN(n418) );
  NAND2_X1 U549 ( .A1(n642), .A2(n585), .ZN(n586) );
  NAND2_X1 U550 ( .A1(n420), .A2(n467), .ZN(n466) );
  NOR2_X1 U551 ( .A1(n653), .A2(KEYINPUT65), .ZN(n420) );
  NAND2_X1 U552 ( .A1(n424), .A2(n583), .ZN(n421) );
  XNOR2_X2 U553 ( .A(n422), .B(n560), .ZN(n779) );
  XNOR2_X1 U554 ( .A(n579), .B(n423), .ZN(n426) );
  XNOR2_X1 U555 ( .A(n643), .B(n644), .ZN(n645) );
  NAND2_X1 U556 ( .A1(n564), .A2(n463), .ZN(n471) );
  XNOR2_X1 U557 ( .A(n561), .B(KEYINPUT108), .ZN(n564) );
  NAND2_X1 U558 ( .A1(n468), .A2(n466), .ZN(n431) );
  XNOR2_X1 U559 ( .A(n432), .B(n646), .ZN(G57) );
  NOR2_X2 U560 ( .A1(n645), .A2(n751), .ZN(n432) );
  NOR2_X2 U561 ( .A1(n598), .A2(n530), .ZN(n462) );
  INV_X1 U562 ( .A(n672), .ZN(n443) );
  XNOR2_X1 U563 ( .A(n433), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U564 ( .A1(n743), .A2(n751), .ZN(n433) );
  XNOR2_X1 U565 ( .A(n434), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U566 ( .A1(n733), .A2(n751), .ZN(n434) );
  NOR2_X1 U567 ( .A1(n616), .A2(n436), .ZN(n435) );
  NOR2_X1 U568 ( .A1(n749), .A2(G902), .ZN(n437) );
  NAND2_X1 U569 ( .A1(n438), .A2(n767), .ZN(n444) );
  XNOR2_X1 U570 ( .A(n586), .B(n439), .ZN(n438) );
  NAND2_X1 U571 ( .A1(n705), .A2(n704), .ZN(n701) );
  NOR2_X2 U572 ( .A1(n780), .A2(KEYINPUT44), .ZN(n565) );
  XNOR2_X2 U573 ( .A(n449), .B(KEYINPUT35), .ZN(n780) );
  NAND2_X1 U574 ( .A1(n450), .A2(n367), .ZN(n449) );
  NAND2_X1 U575 ( .A1(n690), .A2(KEYINPUT33), .ZN(n457) );
  NOR2_X1 U576 ( .A1(n690), .A2(n689), .ZN(n569) );
  INV_X1 U577 ( .A(n689), .ZN(n456) );
  INV_X1 U578 ( .A(KEYINPUT6), .ZN(n459) );
  XNOR2_X1 U579 ( .A(n557), .B(KEYINPUT105), .ZN(n620) );
  NAND2_X1 U580 ( .A1(n461), .A2(n460), .ZN(n558) );
  NAND2_X1 U581 ( .A1(n779), .A2(n472), .ZN(n469) );
  NOR2_X1 U582 ( .A1(n779), .A2(n653), .ZN(n567) );
  INV_X1 U583 ( .A(n779), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n512), .B(n487), .ZN(n488) );
  XOR2_X1 U585 ( .A(KEYINPUT79), .B(n628), .Z(n478) );
  XNOR2_X1 U586 ( .A(KEYINPUT59), .B(KEYINPUT91), .ZN(n479) );
  NOR2_X1 U587 ( .A1(n478), .A2(n632), .ZN(n633) );
  XNOR2_X1 U588 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U589 ( .A(n620), .ZN(n707) );
  XNOR2_X1 U590 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U591 ( .A(KEYINPUT30), .ZN(n613) );
  XNOR2_X1 U592 ( .A(n483), .B(n482), .ZN(n484) );
  NOR2_X1 U593 ( .A1(n597), .A2(n689), .ZN(n614) );
  INV_X1 U594 ( .A(KEYINPUT40), .ZN(n618) );
  XNOR2_X1 U595 ( .A(KEYINPUT63), .B(KEYINPUT89), .ZN(n646) );
  XOR2_X1 U596 ( .A(KEYINPUT77), .B(n481), .Z(n540) );
  NAND2_X1 U597 ( .A1(G210), .A2(n540), .ZN(n483) );
  XOR2_X1 U598 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n482) );
  INV_X1 U599 ( .A(n518), .ZN(n585) );
  NAND2_X1 U600 ( .A1(G227), .A2(n768), .ZN(n486) );
  NOR2_X1 U601 ( .A1(G902), .A2(n734), .ZN(n489) );
  XOR2_X1 U602 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n492) );
  NAND2_X1 U603 ( .A1(n518), .A2(G234), .ZN(n490) );
  XNOR2_X1 U604 ( .A(n490), .B(KEYINPUT20), .ZN(n503) );
  NAND2_X1 U605 ( .A1(n503), .A2(G221), .ZN(n491) );
  XNOR2_X1 U606 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U607 ( .A(KEYINPUT94), .B(n493), .ZN(n686) );
  XOR2_X1 U608 ( .A(G146), .B(G125), .Z(n513) );
  XOR2_X1 U609 ( .A(G110), .B(G128), .Z(n496) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U611 ( .A(n766), .B(n497), .ZN(n502) );
  XOR2_X1 U612 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n500) );
  NAND2_X1 U613 ( .A1(G234), .A2(n768), .ZN(n498) );
  XOR2_X1 U614 ( .A(KEYINPUT8), .B(n498), .Z(n548) );
  NAND2_X1 U615 ( .A1(G221), .A2(n548), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n502), .B(n501), .ZN(n749) );
  NAND2_X1 U618 ( .A1(n503), .A2(G217), .ZN(n505) );
  OR2_X1 U619 ( .A1(n686), .A2(n685), .ZN(n689) );
  XNOR2_X1 U620 ( .A(G472), .B(KEYINPUT97), .ZN(n508) );
  XOR2_X1 U621 ( .A(n513), .B(KEYINPUT17), .Z(n515) );
  NAND2_X1 U622 ( .A1(G224), .A2(n768), .ZN(n514) );
  OR2_X1 U623 ( .A1(G237), .A2(G902), .ZN(n521) );
  NAND2_X1 U624 ( .A1(n521), .A2(G210), .ZN(n519) );
  NAND2_X1 U625 ( .A1(G214), .A2(n521), .ZN(n704) );
  INV_X1 U626 ( .A(n704), .ZN(n602) );
  NAND2_X1 U627 ( .A1(n768), .A2(G952), .ZN(n587) );
  NAND2_X1 U628 ( .A1(G953), .A2(G902), .ZN(n588) );
  OR2_X1 U629 ( .A1(n588), .A2(G898), .ZN(n526) );
  NAND2_X1 U630 ( .A1(n587), .A2(n526), .ZN(n524) );
  XNOR2_X1 U631 ( .A(KEYINPUT14), .B(n523), .ZN(n591) );
  NAND2_X1 U632 ( .A1(n524), .A2(n591), .ZN(n525) );
  NAND2_X1 U633 ( .A1(n525), .A2(KEYINPUT92), .ZN(n529) );
  NOR2_X1 U634 ( .A1(KEYINPUT92), .A2(n526), .ZN(n527) );
  NAND2_X1 U635 ( .A1(n527), .A2(n591), .ZN(n528) );
  NAND2_X1 U636 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U637 ( .A(n531), .B(n766), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n537) );
  XNOR2_X1 U639 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U640 ( .A(n537), .B(n536), .Z(n538) );
  NOR2_X1 U641 ( .A1(G902), .A2(n740), .ZN(n543) );
  XNOR2_X1 U642 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n541) );
  XNOR2_X1 U643 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U644 ( .A(n547), .B(n546), .Z(n550) );
  NAND2_X1 U645 ( .A1(G217), .A2(n548), .ZN(n549) );
  XNOR2_X1 U646 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U647 ( .A(G122), .B(KEYINPUT7), .Z(n551) );
  XNOR2_X1 U648 ( .A(n552), .B(n551), .ZN(n745) );
  NOR2_X1 U649 ( .A1(G902), .A2(n745), .ZN(n553) );
  XNOR2_X1 U650 ( .A(G478), .B(n553), .ZN(n574) );
  INV_X1 U651 ( .A(n574), .ZN(n556) );
  NAND2_X1 U652 ( .A1(n573), .A2(n556), .ZN(n554) );
  XOR2_X1 U653 ( .A(KEYINPUT90), .B(n690), .Z(n610) );
  NAND2_X1 U654 ( .A1(n685), .A2(n610), .ZN(n555) );
  XNOR2_X1 U655 ( .A(KEYINPUT107), .B(n555), .ZN(n559) );
  INV_X1 U656 ( .A(KEYINPUT32), .ZN(n560) );
  INV_X1 U657 ( .A(n693), .ZN(n562) );
  AND2_X1 U658 ( .A1(n685), .A2(n562), .ZN(n563) );
  NAND2_X1 U659 ( .A1(n565), .A2(n567), .ZN(n568) );
  INV_X1 U660 ( .A(KEYINPUT44), .ZN(n566) );
  NAND2_X1 U661 ( .A1(n780), .A2(KEYINPUT44), .ZN(n578) );
  NAND2_X1 U662 ( .A1(n693), .A2(n569), .ZN(n698) );
  XNOR2_X1 U663 ( .A(n570), .B(KEYINPUT31), .ZN(n663) );
  NOR2_X1 U664 ( .A1(n693), .A2(n571), .ZN(n572) );
  NAND2_X1 U665 ( .A1(n614), .A2(n572), .ZN(n648) );
  NAND2_X1 U666 ( .A1(n663), .A2(n648), .ZN(n576) );
  NAND2_X1 U667 ( .A1(n574), .A2(n573), .ZN(n661) );
  OR2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n664) );
  XNOR2_X1 U669 ( .A(KEYINPUT102), .B(n664), .ZN(n634) );
  NAND2_X1 U670 ( .A1(n661), .A2(n634), .ZN(n575) );
  XOR2_X1 U671 ( .A(n575), .B(KEYINPUT103), .Z(n625) );
  NAND2_X1 U672 ( .A1(n576), .A2(n625), .ZN(n577) );
  NAND2_X1 U673 ( .A1(n578), .A2(n577), .ZN(n582) );
  INV_X1 U674 ( .A(n777), .ZN(n581) );
  INV_X1 U675 ( .A(n686), .ZN(n593) );
  INV_X1 U676 ( .A(n587), .ZN(n590) );
  NOR2_X1 U677 ( .A1(G900), .A2(n588), .ZN(n589) );
  NOR2_X1 U678 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U679 ( .A(n591), .ZN(n716) );
  NOR2_X1 U680 ( .A1(n592), .A2(n716), .ZN(n615) );
  NAND2_X1 U681 ( .A1(n593), .A2(n615), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n685), .A2(n693), .ZN(n594) );
  NOR2_X1 U683 ( .A1(n601), .A2(n594), .ZN(n595) );
  XOR2_X1 U684 ( .A(KEYINPUT28), .B(n595), .Z(n596) );
  NOR2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n621) );
  INV_X1 U686 ( .A(n598), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n621), .A2(n599), .ZN(n659) );
  NAND2_X1 U688 ( .A1(n659), .A2(KEYINPUT47), .ZN(n600) );
  XNOR2_X1 U689 ( .A(n600), .B(KEYINPUT80), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT36), .B(KEYINPUT88), .Z(n608) );
  NOR2_X1 U691 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U692 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n661), .A2(n605), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n685), .A2(n606), .ZN(n637) );
  NOR2_X1 U695 ( .A1(n441), .A2(n637), .ZN(n607) );
  XOR2_X1 U696 ( .A(n608), .B(n607), .Z(n609) );
  NAND2_X1 U697 ( .A1(n610), .A2(n609), .ZN(n667) );
  XOR2_X1 U698 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n612) );
  XNOR2_X1 U699 ( .A(KEYINPUT86), .B(n612), .ZN(n623) );
  XNOR2_X1 U700 ( .A(KEYINPUT38), .B(n441), .ZN(n705) );
  XNOR2_X1 U701 ( .A(n617), .B(n375), .ZN(n635) );
  NOR2_X1 U702 ( .A1(n635), .A2(n661), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n441), .A2(n624), .ZN(n658) );
  XNOR2_X1 U704 ( .A(n658), .B(KEYINPUT81), .ZN(n627) );
  INV_X1 U705 ( .A(n625), .ZN(n702) );
  NAND2_X1 U706 ( .A1(n702), .A2(KEYINPUT47), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U708 ( .A1(KEYINPUT47), .A2(n702), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n629), .B(KEYINPUT75), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n659), .A2(n630), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n631), .B(KEYINPUT74), .ZN(n632) );
  NOR2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n668) );
  XOR2_X1 U713 ( .A(n637), .B(KEYINPUT110), .Z(n638) );
  NAND2_X1 U714 ( .A1(n638), .A2(n690), .ZN(n639) );
  XNOR2_X1 U715 ( .A(n639), .B(KEYINPUT43), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n641), .A2(n441), .ZN(n669) );
  NAND2_X1 U717 ( .A1(n747), .A2(G472), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n661), .A2(n648), .ZN(n647) );
  XOR2_X1 U719 ( .A(G104), .B(n647), .Z(G6) );
  NOR2_X1 U720 ( .A1(n648), .A2(n664), .ZN(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n650) );
  XNOR2_X1 U722 ( .A(G107), .B(KEYINPUT113), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(G9) );
  XOR2_X1 U725 ( .A(G110), .B(n653), .Z(G12) );
  NOR2_X1 U726 ( .A1(n659), .A2(n664), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n655) );
  XNOR2_X1 U728 ( .A(G128), .B(KEYINPUT115), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(G30) );
  XOR2_X1 U731 ( .A(G143), .B(n658), .Z(G45) );
  NOR2_X1 U732 ( .A1(n661), .A2(n659), .ZN(n660) );
  XOR2_X1 U733 ( .A(G146), .B(n660), .Z(G48) );
  NOR2_X1 U734 ( .A1(n661), .A2(n663), .ZN(n662) );
  XOR2_X1 U735 ( .A(G113), .B(n662), .Z(G15) );
  NOR2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U737 ( .A(G116), .B(n665), .Z(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(G27) );
  XOR2_X1 U740 ( .A(G134), .B(n668), .Z(G36) );
  XNOR2_X1 U741 ( .A(G140), .B(KEYINPUT116), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(G42) );
  XOR2_X1 U743 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n727) );
  INV_X1 U744 ( .A(KEYINPUT82), .ZN(n677) );
  AND2_X1 U745 ( .A1(n677), .A2(n752), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n684) );
  NAND2_X1 U747 ( .A1(n767), .A2(KEYINPUT83), .ZN(n676) );
  OR2_X1 U748 ( .A1(n677), .A2(KEYINPUT83), .ZN(n674) );
  NAND2_X1 U749 ( .A1(KEYINPUT2), .A2(n674), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n682) );
  NOR2_X1 U751 ( .A1(n767), .A2(KEYINPUT83), .ZN(n679) );
  NOR2_X1 U752 ( .A1(n752), .A2(n677), .ZN(n678) );
  NOR2_X1 U753 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U754 ( .A1(KEYINPUT2), .A2(n680), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n719) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(KEYINPUT117), .ZN(n688) );
  XNOR2_X1 U759 ( .A(KEYINPUT49), .B(n688), .ZN(n696) );
  XOR2_X1 U760 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n692) );
  NAND2_X1 U761 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U766 ( .A(KEYINPUT51), .B(n699), .Z(n700) );
  NAND2_X1 U767 ( .A1(n721), .A2(n700), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT120), .B(n703), .Z(n710) );
  NOR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U771 ( .A(KEYINPUT119), .B(n706), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U774 ( .A1(n720), .A2(n711), .ZN(n712) );
  NAND2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U776 ( .A(KEYINPUT52), .B(n714), .Z(n715) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n717), .A2(G952), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(KEYINPUT121), .B(n722), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U783 ( .A1(n725), .A2(n768), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n727), .B(n726), .ZN(G75) );
  NAND2_X1 U785 ( .A1(n747), .A2(G210), .ZN(n732) );
  INV_X1 U786 ( .A(n728), .ZN(n730) );
  XOR2_X1 U787 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n729) );
  XNOR2_X1 U788 ( .A(n732), .B(n731), .ZN(n733) );
  XOR2_X1 U789 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n736) );
  XNOR2_X1 U790 ( .A(n734), .B(KEYINPUT123), .ZN(n735) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n738) );
  NAND2_X1 U792 ( .A1(n747), .A2(G469), .ZN(n737) );
  XOR2_X1 U793 ( .A(n738), .B(n737), .Z(n739) );
  NOR2_X1 U794 ( .A1(n751), .A2(n739), .ZN(G54) );
  NAND2_X1 U795 ( .A1(n747), .A2(G475), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U797 ( .A1(G478), .A2(n360), .ZN(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n751), .A2(n746), .ZN(G63) );
  NAND2_X1 U800 ( .A1(G217), .A2(n360), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n751), .A2(n750), .ZN(G66) );
  NAND2_X1 U803 ( .A1(n768), .A2(n752), .ZN(n756) );
  NAND2_X1 U804 ( .A1(G953), .A2(G224), .ZN(n753) );
  XNOR2_X1 U805 ( .A(KEYINPUT61), .B(n753), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n754), .A2(G898), .ZN(n755) );
  NAND2_X1 U807 ( .A1(n756), .A2(n755), .ZN(n763) );
  NOR2_X1 U808 ( .A1(G898), .A2(n768), .ZN(n761) );
  XOR2_X1 U809 ( .A(n361), .B(G101), .Z(n758) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(G69) );
  XOR2_X1 U813 ( .A(KEYINPUT4), .B(n764), .Z(n765) );
  XOR2_X1 U814 ( .A(n766), .B(n765), .Z(n770) );
  XOR2_X1 U815 ( .A(n770), .B(n767), .Z(n769) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(n776) );
  XNOR2_X1 U817 ( .A(n770), .B(KEYINPUT124), .ZN(n771) );
  XNOR2_X1 U818 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U819 ( .A1(G900), .A2(n772), .ZN(n773) );
  XOR2_X1 U820 ( .A(KEYINPUT125), .B(n773), .Z(n774) );
  NAND2_X1 U821 ( .A1(G953), .A2(n774), .ZN(n775) );
  NAND2_X1 U822 ( .A1(n776), .A2(n775), .ZN(G72) );
  XNOR2_X1 U823 ( .A(n777), .B(G101), .ZN(n778) );
  XNOR2_X1 U824 ( .A(n778), .B(KEYINPUT112), .ZN(G3) );
  XOR2_X1 U825 ( .A(G119), .B(n779), .Z(G21) );
  XOR2_X1 U826 ( .A(n780), .B(G122), .Z(n781) );
  XNOR2_X1 U827 ( .A(KEYINPUT126), .B(n781), .ZN(G24) );
  XNOR2_X1 U828 ( .A(G137), .B(n782), .ZN(G39) );
endmodule

