

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809;

  AND2_X1 U379 ( .A1(n655), .A2(n532), .ZN(n446) );
  OR2_X2 U380 ( .A1(n666), .A2(n732), .ZN(n579) );
  NOR2_X2 U381 ( .A1(n642), .A2(n636), .ZN(n492) );
  XNOR2_X2 U382 ( .A(n537), .B(G131), .ZN(n581) );
  XNOR2_X2 U383 ( .A(G146), .B(KEYINPUT68), .ZN(n537) );
  XNOR2_X2 U384 ( .A(n582), .B(G119), .ZN(n489) );
  XNOR2_X2 U385 ( .A(KEYINPUT3), .B(KEYINPUT71), .ZN(n582) );
  XNOR2_X2 U386 ( .A(n442), .B(n517), .ZN(n694) );
  XNOR2_X2 U387 ( .A(n391), .B(n791), .ZN(n442) );
  XNOR2_X2 U388 ( .A(G107), .B(G104), .ZN(n528) );
  NOR2_X2 U389 ( .A1(G902), .A2(n767), .ZN(n595) );
  INV_X1 U390 ( .A(G953), .ZN(n797) );
  NOR2_X2 U391 ( .A1(G953), .A2(G237), .ZN(n540) );
  XNOR2_X1 U392 ( .A(n445), .B(n656), .ZN(n658) );
  XNOR2_X1 U393 ( .A(n491), .B(KEYINPUT40), .ZN(n806) );
  NAND2_X1 U394 ( .A1(n658), .A2(n529), .ZN(n401) );
  AND2_X1 U395 ( .A1(n462), .A2(KEYINPUT66), .ZN(n437) );
  NAND2_X1 U396 ( .A1(n369), .A2(n425), .ZN(n424) );
  AND2_X1 U397 ( .A1(n511), .A2(KEYINPUT32), .ZN(n409) );
  AND2_X1 U398 ( .A1(n516), .A2(n515), .ZN(n514) );
  NOR2_X1 U399 ( .A1(n753), .A2(KEYINPUT47), .ZN(n648) );
  AND2_X1 U400 ( .A1(n627), .A2(n626), .ZN(n644) );
  XNOR2_X1 U401 ( .A(n459), .B(n633), .ZN(n738) );
  XNOR2_X1 U402 ( .A(n573), .B(KEYINPUT25), .ZN(n574) );
  NAND2_X1 U403 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U404 ( .A(n495), .B(KEYINPUT10), .ZN(n564) );
  XNOR2_X1 U405 ( .A(G125), .B(G140), .ZN(n495) );
  INV_X1 U406 ( .A(KEYINPUT33), .ZN(n433) );
  INV_X1 U407 ( .A(n634), .ZN(n359) );
  NOR2_X1 U408 ( .A1(n360), .A2(n738), .ZN(n635) );
  NAND2_X1 U409 ( .A1(n626), .A2(n359), .ZN(n360) );
  NOR2_X1 U410 ( .A1(n779), .A2(G902), .ZN(n575) );
  BUF_X1 U411 ( .A(n806), .Z(n361) );
  BUF_X1 U412 ( .A(n796), .Z(n362) );
  BUF_X1 U413 ( .A(n786), .Z(n363) );
  XNOR2_X1 U414 ( .A(n526), .B(KEYINPUT19), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n599), .B(n443), .ZN(n786) );
  NAND2_X2 U416 ( .A1(n497), .A2(n508), .ZN(n526) );
  BUF_X1 U417 ( .A(n671), .Z(n365) );
  XNOR2_X1 U418 ( .A(n494), .B(n493), .ZN(n563) );
  INV_X1 U419 ( .A(KEYINPUT8), .ZN(n493) );
  NAND2_X1 U420 ( .A1(n507), .A2(n606), .ZN(n506) );
  NAND2_X1 U421 ( .A1(n609), .A2(n685), .ZN(n509) );
  AND2_X1 U422 ( .A1(n485), .A2(n663), .ZN(n484) );
  INV_X1 U423 ( .A(KEYINPUT36), .ZN(n408) );
  AND2_X1 U424 ( .A1(n623), .A2(n482), .ZN(n498) );
  XNOR2_X1 U425 ( .A(n805), .B(KEYINPUT84), .ZN(n451) );
  INV_X1 U426 ( .A(G237), .ZN(n589) );
  XNOR2_X1 U427 ( .A(n545), .B(n368), .ZN(n518) );
  INV_X1 U428 ( .A(KEYINPUT6), .ZN(n463) );
  XNOR2_X1 U429 ( .A(n584), .B(n585), .ZN(n490) );
  XNOR2_X1 U430 ( .A(G116), .B(G113), .ZN(n488) );
  XNOR2_X1 U431 ( .A(n449), .B(n570), .ZN(n779) );
  XNOR2_X1 U432 ( .A(n793), .B(n450), .ZN(n449) );
  XNOR2_X1 U433 ( .A(n555), .B(KEYINPUT9), .ZN(n522) );
  XNOR2_X1 U434 ( .A(G116), .B(G122), .ZN(n555) );
  INV_X1 U435 ( .A(KEYINPUT65), .ZN(n477) );
  XNOR2_X1 U436 ( .A(n392), .B(n391), .ZN(n702) );
  XNOR2_X1 U437 ( .A(n625), .B(n480), .ZN(n627) );
  XNOR2_X1 U438 ( .A(n481), .B(KEYINPUT28), .ZN(n480) );
  AND2_X1 U439 ( .A1(n419), .A2(n417), .ZN(n422) );
  AND2_X1 U440 ( .A1(n591), .A2(n376), .ZN(n406) );
  INV_X1 U441 ( .A(KEYINPUT32), .ZN(n461) );
  NAND2_X1 U442 ( .A1(n414), .A2(KEYINPUT32), .ZN(n413) );
  INV_X1 U443 ( .A(n498), .ZN(n414) );
  XNOR2_X1 U444 ( .A(n557), .B(G478), .ZN(n645) );
  NOR2_X1 U445 ( .A1(n774), .A2(G902), .ZN(n557) );
  NAND2_X1 U446 ( .A1(n646), .A2(n645), .ZN(n638) );
  INV_X1 U447 ( .A(KEYINPUT1), .ZN(n435) );
  XNOR2_X1 U448 ( .A(n504), .B(n502), .ZN(n594) );
  XNOR2_X1 U449 ( .A(n592), .B(n503), .ZN(n502) );
  XNOR2_X1 U450 ( .A(n394), .B(KEYINPUT83), .ZN(n393) );
  INV_X1 U451 ( .A(KEYINPUT90), .ZN(n441) );
  XNOR2_X1 U452 ( .A(G113), .B(G104), .ZN(n535) );
  INV_X1 U453 ( .A(G902), .ZN(n590) );
  OR2_X1 U454 ( .A1(n752), .A2(n732), .ZN(n620) );
  INV_X1 U455 ( .A(KEYINPUT44), .ZN(n440) );
  XNOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT79), .ZN(n567) );
  XNOR2_X1 U457 ( .A(n564), .B(n593), .ZN(n793) );
  NAND2_X1 U458 ( .A1(n563), .A2(G221), .ZN(n450) );
  XNOR2_X1 U459 ( .A(G119), .B(G128), .ZN(n565) );
  XNOR2_X1 U460 ( .A(n478), .B(n536), .ZN(n539) );
  XOR2_X1 U461 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n536) );
  XNOR2_X1 U462 ( .A(n535), .B(n479), .ZN(n478) );
  INV_X1 U463 ( .A(G122), .ZN(n479) );
  NOR2_X1 U464 ( .A1(n395), .A2(n396), .ZN(n687) );
  XOR2_X1 U465 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n601) );
  XNOR2_X1 U466 ( .A(G146), .B(G125), .ZN(n600) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n558) );
  INV_X1 U468 ( .A(KEYINPUT107), .ZN(n481) );
  NAND2_X1 U469 ( .A1(n423), .A2(n749), .ZN(n421) );
  OR2_X1 U470 ( .A1(n750), .A2(n423), .ZN(n419) );
  OR2_X1 U471 ( .A1(n752), .A2(n611), .ZN(n418) );
  NOR2_X1 U472 ( .A1(n620), .A2(n622), .ZN(n512) );
  INV_X1 U473 ( .A(KEYINPUT30), .ZN(n468) );
  XNOR2_X1 U474 ( .A(n526), .B(KEYINPUT19), .ZN(n643) );
  XOR2_X1 U475 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n572) );
  INV_X1 U476 ( .A(KEYINPUT80), .ZN(n503) );
  INV_X1 U477 ( .A(KEYINPUT39), .ZN(n637) );
  AND2_X1 U478 ( .A1(n484), .A2(KEYINPUT35), .ZN(n431) );
  XNOR2_X1 U479 ( .A(n586), .B(G137), .ZN(n517) );
  XNOR2_X1 U480 ( .A(n490), .B(n388), .ZN(n586) );
  XNOR2_X1 U481 ( .A(n496), .B(n598), .ZN(n599) );
  XNOR2_X1 U482 ( .A(n521), .B(n519), .ZN(n774) );
  XNOR2_X1 U483 ( .A(n554), .B(n520), .ZN(n519) );
  XNOR2_X1 U484 ( .A(n556), .B(n522), .ZN(n521) );
  XNOR2_X1 U485 ( .A(n531), .B(n629), .ZN(n808) );
  NAND2_X1 U486 ( .A1(n651), .A2(n375), .ZN(n405) );
  AND2_X1 U487 ( .A1(n498), .A2(n461), .ZN(n460) );
  XNOR2_X1 U488 ( .A(n453), .B(n452), .ZN(n805) );
  NAND2_X1 U489 ( .A1(n670), .A2(n482), .ZN(n681) );
  INV_X1 U490 ( .A(KEYINPUT124), .ZN(n472) );
  INV_X1 U491 ( .A(KEYINPUT60), .ZN(n469) );
  XNOR2_X1 U492 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U493 ( .A1(n765), .A2(G953), .ZN(n471) );
  AND2_X1 U494 ( .A1(n438), .A2(n378), .ZN(n366) );
  INV_X1 U495 ( .A(KEYINPUT35), .ZN(n664) );
  NOR2_X1 U496 ( .A1(n486), .A2(n675), .ZN(n367) );
  XOR2_X1 U497 ( .A(KEYINPUT13), .B(G475), .Z(n368) );
  AND2_X1 U498 ( .A1(n432), .A2(n431), .ZN(n369) );
  XOR2_X1 U499 ( .A(KEYINPUT120), .B(n729), .Z(n370) );
  AND2_X1 U500 ( .A1(n518), .A2(n645), .ZN(n371) );
  XOR2_X1 U501 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n372) );
  XOR2_X1 U502 ( .A(n693), .B(n692), .Z(n373) );
  AND2_X1 U503 ( .A1(n530), .A2(n691), .ZN(n374) );
  OR2_X1 U504 ( .A1(n407), .A2(n408), .ZN(n375) );
  AND2_X1 U505 ( .A1(n407), .A2(n408), .ZN(n376) );
  AND2_X1 U506 ( .A1(n626), .A2(n500), .ZN(n377) );
  AND2_X1 U507 ( .A1(n682), .A2(n708), .ZN(n378) );
  NOR2_X1 U508 ( .A1(n752), .A2(n421), .ZN(n379) );
  NOR2_X1 U509 ( .A1(n763), .A2(n370), .ZN(n380) );
  XOR2_X1 U510 ( .A(KEYINPUT70), .B(G469), .Z(n381) );
  XNOR2_X1 U511 ( .A(KEYINPUT46), .B(KEYINPUT89), .ZN(n382) );
  XOR2_X1 U512 ( .A(n628), .B(KEYINPUT41), .Z(n383) );
  INV_X1 U513 ( .A(KEYINPUT34), .ZN(n524) );
  XNOR2_X1 U514 ( .A(n779), .B(KEYINPUT123), .ZN(n384) );
  INV_X1 U515 ( .A(n606), .ZN(n685) );
  XNOR2_X1 U516 ( .A(G902), .B(KEYINPUT15), .ZN(n606) );
  NOR2_X1 U517 ( .A1(KEYINPUT85), .A2(n606), .ZN(n385) );
  AND2_X1 U518 ( .A1(n697), .A2(G953), .ZN(n781) );
  INV_X1 U519 ( .A(n781), .ZN(n474) );
  XNOR2_X2 U520 ( .A(KEYINPUT103), .B(n647), .ZN(n753) );
  XNOR2_X1 U521 ( .A(n771), .B(KEYINPUT59), .ZN(n534) );
  AND2_X1 U522 ( .A1(n658), .A2(n657), .ZN(n530) );
  NOR2_X1 U523 ( .A1(G902), .A2(n771), .ZN(n545) );
  NAND2_X1 U524 ( .A1(n426), .A2(n424), .ZN(n386) );
  NAND2_X1 U525 ( .A1(n426), .A2(n424), .ZN(n462) );
  AND2_X1 U526 ( .A1(n672), .A2(n524), .ZN(n487) );
  AND2_X2 U527 ( .A1(n476), .A2(n373), .ZN(n387) );
  XNOR2_X1 U528 ( .A(n489), .B(n488), .ZN(n388) );
  XNOR2_X2 U529 ( .A(n465), .B(n477), .ZN(n476) );
  XNOR2_X1 U530 ( .A(n489), .B(n488), .ZN(n443) );
  AND2_X1 U531 ( .A1(n454), .A2(n451), .ZN(n655) );
  XNOR2_X1 U532 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U533 ( .A1(n649), .A2(n611), .ZN(n407) );
  XNOR2_X1 U534 ( .A(n649), .B(KEYINPUT38), .ZN(n750) );
  OR2_X2 U535 ( .A1(n702), .A2(n506), .ZN(n505) );
  XNOR2_X1 U536 ( .A(n630), .B(n463), .ZN(n464) );
  INV_X1 U537 ( .A(n738), .ZN(n500) );
  NAND2_X1 U538 ( .A1(n666), .A2(n632), .ZN(n459) );
  XNOR2_X1 U539 ( .A(n455), .B(KEYINPUT74), .ZN(n454) );
  NAND2_X1 U540 ( .A1(n475), .A2(n474), .ZN(n473) );
  XNOR2_X1 U541 ( .A(n780), .B(n384), .ZN(n475) );
  BUF_X1 U542 ( .A(n750), .Z(n416) );
  NOR2_X1 U543 ( .A1(n683), .A2(KEYINPUT2), .ZN(n394) );
  NAND2_X1 U544 ( .A1(n460), .A2(n411), .ZN(n410) );
  NAND2_X1 U545 ( .A1(n672), .A2(n512), .ZN(n389) );
  NAND2_X1 U546 ( .A1(n513), .A2(n512), .ZN(n511) );
  INV_X1 U547 ( .A(n580), .ZN(n520) );
  XNOR2_X1 U548 ( .A(n448), .B(n441), .ZN(n390) );
  XNOR2_X1 U549 ( .A(n448), .B(n441), .ZN(n397) );
  XNOR2_X1 U550 ( .A(n786), .B(n605), .ZN(n392) );
  XNOR2_X2 U551 ( .A(n795), .B(G101), .ZN(n391) );
  NAND2_X1 U552 ( .A1(n702), .A2(n609), .ZN(n510) );
  NAND2_X1 U553 ( .A1(n393), .A2(n373), .ZN(n466) );
  INV_X1 U554 ( .A(n398), .ZN(n395) );
  NAND2_X1 U555 ( .A1(n796), .A2(n385), .ZN(n396) );
  AND2_X2 U556 ( .A1(n796), .A2(n398), .ZN(n683) );
  NAND2_X1 U557 ( .A1(n397), .A2(n437), .ZN(n402) );
  NAND2_X1 U558 ( .A1(n439), .A2(n390), .ZN(n438) );
  NAND2_X1 U559 ( .A1(n398), .A2(n374), .ZN(n693) );
  NAND2_X1 U560 ( .A1(n398), .A2(n797), .ZN(n785) );
  XNOR2_X2 U561 ( .A(n399), .B(KEYINPUT45), .ZN(n398) );
  NAND2_X1 U562 ( .A1(n400), .A2(n366), .ZN(n399) );
  XNOR2_X1 U563 ( .A(n402), .B(n440), .ZN(n400) );
  XNOR2_X2 U564 ( .A(n401), .B(n662), .ZN(n796) );
  XNOR2_X1 U565 ( .A(n631), .B(n468), .ZN(n467) );
  NAND2_X1 U566 ( .A1(n404), .A2(n403), .ZN(n728) );
  OR2_X1 U567 ( .A1(n591), .A2(n408), .ZN(n403) );
  NOR2_X1 U568 ( .A1(n406), .A2(n405), .ZN(n404) );
  NAND2_X1 U569 ( .A1(n591), .A2(n749), .ZN(n650) );
  NAND2_X1 U570 ( .A1(n409), .A2(n514), .ZN(n415) );
  NAND2_X2 U571 ( .A1(n412), .A2(n410), .ZN(n671) );
  NAND2_X1 U572 ( .A1(n514), .A2(n389), .ZN(n411) );
  AND2_X2 U573 ( .A1(n415), .A2(n413), .ZN(n412) );
  XNOR2_X2 U574 ( .A(n595), .B(n381), .ZN(n626) );
  NAND2_X1 U575 ( .A1(n418), .A2(n383), .ZN(n417) );
  NAND2_X1 U576 ( .A1(n416), .A2(n749), .ZN(n444) );
  NAND2_X1 U577 ( .A1(n422), .A2(n420), .ZN(n747) );
  NAND2_X1 U578 ( .A1(n416), .A2(n379), .ZN(n420) );
  INV_X1 U579 ( .A(n383), .ZN(n423) );
  NAND2_X1 U580 ( .A1(n487), .A2(n434), .ZN(n432) );
  NAND2_X1 U581 ( .A1(n483), .A2(KEYINPUT34), .ZN(n425) );
  AND2_X2 U582 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U583 ( .A1(n483), .A2(n430), .ZN(n427) );
  NAND2_X1 U584 ( .A1(n429), .A2(n664), .ZN(n428) );
  NAND2_X1 U585 ( .A1(n432), .A2(n484), .ZN(n429) );
  NOR2_X1 U586 ( .A1(n524), .A2(KEYINPUT35), .ZN(n430) );
  INV_X1 U587 ( .A(n434), .ZN(n483) );
  XNOR2_X2 U588 ( .A(n525), .B(n433), .ZN(n434) );
  NAND2_X1 U589 ( .A1(n757), .A2(n434), .ZN(n758) );
  XNOR2_X2 U590 ( .A(n626), .B(n435), .ZN(n737) );
  OR2_X1 U591 ( .A1(n483), .A2(n436), .ZN(n729) );
  INV_X1 U592 ( .A(n747), .ZN(n436) );
  OR2_X2 U593 ( .A1(n724), .A2(n722), .ZN(n647) );
  AND2_X2 U594 ( .A1(n476), .A2(n373), .ZN(n778) );
  NOR2_X1 U595 ( .A1(n386), .A2(KEYINPUT66), .ZN(n439) );
  XNOR2_X1 U596 ( .A(n442), .B(n523), .ZN(n767) );
  NOR2_X1 U597 ( .A1(n753), .A2(n444), .ZN(n754) );
  NAND2_X1 U598 ( .A1(n447), .A2(n446), .ZN(n445) );
  XNOR2_X1 U599 ( .A(n639), .B(n382), .ZN(n447) );
  NAND2_X2 U600 ( .A1(n671), .A2(n716), .ZN(n448) );
  INV_X1 U601 ( .A(KEYINPUT106), .ZN(n452) );
  NOR2_X1 U602 ( .A1(n642), .A2(n641), .ZN(n453) );
  NAND2_X1 U603 ( .A1(n457), .A2(n456), .ZN(n455) );
  INV_X1 U604 ( .A(n652), .ZN(n456) );
  XNOR2_X1 U605 ( .A(n648), .B(n458), .ZN(n457) );
  INV_X1 U606 ( .A(KEYINPUT75), .ZN(n458) );
  NAND2_X1 U607 ( .A1(n514), .A2(n389), .ZN(n670) );
  XNOR2_X1 U608 ( .A(n386), .B(G122), .ZN(G24) );
  NAND2_X1 U609 ( .A1(n464), .A2(n500), .ZN(n499) );
  INV_X1 U610 ( .A(n464), .ZN(n482) );
  NAND2_X1 U611 ( .A1(n464), .A2(n624), .ZN(n588) );
  INV_X1 U612 ( .A(n750), .ZN(n636) );
  NAND2_X1 U613 ( .A1(n676), .A2(KEYINPUT34), .ZN(n485) );
  NAND2_X1 U614 ( .A1(n688), .A2(n689), .ZN(n465) );
  NAND2_X1 U615 ( .A1(n466), .A2(n380), .ZN(n764) );
  NAND2_X2 U616 ( .A1(n508), .A2(n505), .ZN(n649) );
  NAND2_X1 U617 ( .A1(n635), .A2(n467), .ZN(n642) );
  XNOR2_X1 U618 ( .A(n470), .B(n469), .ZN(G60) );
  NAND2_X1 U619 ( .A1(n773), .A2(n474), .ZN(n470) );
  XNOR2_X1 U620 ( .A(n471), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U621 ( .A(n473), .B(n472), .ZN(G66) );
  INV_X1 U622 ( .A(n518), .ZN(n646) );
  INV_X1 U623 ( .A(n672), .ZN(n486) );
  NAND2_X1 U624 ( .A1(n659), .A2(n722), .ZN(n491) );
  XNOR2_X1 U625 ( .A(n492), .B(n637), .ZN(n659) );
  NAND2_X1 U626 ( .A1(n797), .A2(G234), .ZN(n494) );
  XNOR2_X1 U627 ( .A(n496), .B(n593), .ZN(n504) );
  XNOR2_X2 U628 ( .A(n528), .B(n527), .ZN(n496) );
  AND2_X2 U629 ( .A1(n505), .A2(n749), .ZN(n497) );
  OR2_X1 U630 ( .A1(n737), .A2(n738), .ZN(n501) );
  NOR2_X2 U631 ( .A1(n499), .A2(n737), .ZN(n525) );
  NOR2_X1 U632 ( .A1(n501), .A2(n665), .ZN(n745) );
  INV_X1 U633 ( .A(n609), .ZN(n507) );
  AND2_X2 U634 ( .A1(n510), .A2(n509), .ZN(n508) );
  INV_X1 U635 ( .A(n676), .ZN(n513) );
  NAND2_X1 U636 ( .A1(n620), .A2(n622), .ZN(n515) );
  NAND2_X1 U637 ( .A1(n676), .A2(n622), .ZN(n516) );
  XNOR2_X2 U638 ( .A(n618), .B(n617), .ZN(n676) );
  INV_X1 U639 ( .A(n630), .ZN(n665) );
  NOR2_X1 U640 ( .A1(n645), .A2(n518), .ZN(n663) );
  XNOR2_X1 U641 ( .A(n594), .B(G140), .ZN(n523) );
  NAND2_X1 U642 ( .A1(n643), .A2(n616), .ZN(n618) );
  XNOR2_X2 U643 ( .A(KEYINPUT76), .B(G110), .ZN(n527) );
  AND2_X1 U644 ( .A1(n657), .A2(n661), .ZN(n529) );
  NAND2_X1 U645 ( .A1(n806), .A2(n808), .ZN(n639) );
  NAND2_X1 U646 ( .A1(n644), .A2(n747), .ZN(n531) );
  XNOR2_X1 U647 ( .A(n767), .B(n766), .ZN(n768) );
  AND2_X1 U648 ( .A1(n728), .A2(n654), .ZN(n532) );
  XNOR2_X1 U649 ( .A(G472), .B(KEYINPUT100), .ZN(n533) );
  INV_X1 U650 ( .A(n564), .ZN(n541) );
  INV_X1 U651 ( .A(KEYINPUT108), .ZN(n628) );
  XNOR2_X1 U652 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U653 ( .A(n544), .B(n543), .ZN(n771) );
  XNOR2_X1 U654 ( .A(G143), .B(n581), .ZN(n538) );
  XNOR2_X1 U655 ( .A(n539), .B(n538), .ZN(n544) );
  XOR2_X1 U656 ( .A(KEYINPUT77), .B(n540), .Z(n583) );
  NAND2_X1 U657 ( .A1(G214), .A2(n583), .ZN(n542) );
  INV_X1 U658 ( .A(G128), .ZN(n546) );
  NAND2_X1 U659 ( .A1(n546), .A2(KEYINPUT81), .ZN(n549) );
  INV_X1 U660 ( .A(KEYINPUT81), .ZN(n547) );
  NAND2_X1 U661 ( .A1(n547), .A2(G128), .ZN(n548) );
  XNOR2_X2 U662 ( .A(G143), .B(KEYINPUT64), .ZN(n550) );
  XNOR2_X2 U663 ( .A(n551), .B(n550), .ZN(n580) );
  NAND2_X1 U664 ( .A1(n563), .A2(G217), .ZN(n556) );
  XOR2_X1 U665 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n553) );
  XNOR2_X1 U666 ( .A(G134), .B(G107), .ZN(n552) );
  XNOR2_X1 U667 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U668 ( .A(n558), .B(KEYINPUT14), .ZN(n559) );
  NAND2_X1 U669 ( .A1(G952), .A2(n559), .ZN(n762) );
  NOR2_X1 U670 ( .A1(n762), .A2(G953), .ZN(n613) );
  NAND2_X1 U671 ( .A1(n559), .A2(G902), .ZN(n560) );
  XNOR2_X1 U672 ( .A(n560), .B(KEYINPUT95), .ZN(n612) );
  NAND2_X1 U673 ( .A1(G953), .A2(n612), .ZN(n561) );
  NOR2_X1 U674 ( .A1(G900), .A2(n561), .ZN(n562) );
  NOR2_X1 U675 ( .A1(n613), .A2(n562), .ZN(n634) );
  XOR2_X1 U676 ( .A(G137), .B(KEYINPUT69), .Z(n593) );
  XOR2_X1 U677 ( .A(G110), .B(G146), .Z(n566) );
  XNOR2_X1 U678 ( .A(n566), .B(n565), .ZN(n569) );
  XNOR2_X1 U679 ( .A(n372), .B(n567), .ZN(n568) );
  XOR2_X1 U680 ( .A(n569), .B(n568), .Z(n570) );
  NAND2_X1 U681 ( .A1(G234), .A2(n606), .ZN(n571) );
  XNOR2_X1 U682 ( .A(n572), .B(n571), .ZN(n576) );
  NAND2_X1 U683 ( .A1(G217), .A2(n576), .ZN(n573) );
  XNOR2_X2 U684 ( .A(n575), .B(n574), .ZN(n666) );
  AND2_X1 U685 ( .A1(n576), .A2(G221), .ZN(n578) );
  XNOR2_X1 U686 ( .A(KEYINPUT98), .B(KEYINPUT21), .ZN(n577) );
  XNOR2_X1 U687 ( .A(n578), .B(n577), .ZN(n632) );
  INV_X1 U688 ( .A(n632), .ZN(n732) );
  NOR2_X1 U689 ( .A1(n634), .A2(n579), .ZN(n624) );
  XNOR2_X2 U690 ( .A(n580), .B(KEYINPUT4), .ZN(n795) );
  XNOR2_X1 U691 ( .A(n581), .B(G134), .ZN(n791) );
  NAND2_X1 U692 ( .A1(G210), .A2(n583), .ZN(n584) );
  XOR2_X1 U693 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n585) );
  NAND2_X1 U694 ( .A1(n694), .A2(n590), .ZN(n587) );
  XNOR2_X2 U695 ( .A(n587), .B(n533), .ZN(n630) );
  NOR2_X1 U696 ( .A1(n638), .A2(n588), .ZN(n591) );
  NAND2_X1 U697 ( .A1(n590), .A2(n589), .ZN(n607) );
  NAND2_X1 U698 ( .A1(n607), .A2(G214), .ZN(n749) );
  NAND2_X1 U699 ( .A1(G227), .A2(n797), .ZN(n592) );
  INV_X1 U700 ( .A(n737), .ZN(n651) );
  OR2_X1 U701 ( .A1(n650), .A2(n651), .ZN(n596) );
  XNOR2_X1 U702 ( .A(KEYINPUT43), .B(n596), .ZN(n610) );
  XNOR2_X1 U703 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n597) );
  XNOR2_X1 U704 ( .A(n597), .B(G122), .ZN(n598) );
  XNOR2_X1 U705 ( .A(n601), .B(n600), .ZN(n604) );
  NAND2_X1 U706 ( .A1(n797), .A2(G224), .ZN(n602) );
  XNOR2_X1 U707 ( .A(n602), .B(KEYINPUT93), .ZN(n603) );
  XNOR2_X1 U708 ( .A(n604), .B(n603), .ZN(n605) );
  NAND2_X1 U709 ( .A1(n607), .A2(G210), .ZN(n608) );
  XNOR2_X1 U710 ( .A(n608), .B(KEYINPUT94), .ZN(n609) );
  NAND2_X1 U711 ( .A1(n610), .A2(n649), .ZN(n657) );
  XNOR2_X1 U712 ( .A(n657), .B(G140), .ZN(G42) );
  INV_X1 U713 ( .A(n749), .ZN(n611) );
  NOR2_X1 U714 ( .A1(G898), .A2(n797), .ZN(n787) );
  NAND2_X1 U715 ( .A1(n612), .A2(n787), .ZN(n615) );
  INV_X1 U716 ( .A(n613), .ZN(n614) );
  NAND2_X1 U717 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U718 ( .A(KEYINPUT92), .B(KEYINPUT0), .ZN(n617) );
  INV_X1 U719 ( .A(KEYINPUT104), .ZN(n619) );
  XNOR2_X1 U720 ( .A(n371), .B(n619), .ZN(n752) );
  INV_X1 U721 ( .A(KEYINPUT72), .ZN(n621) );
  XNOR2_X1 U722 ( .A(n621), .B(KEYINPUT22), .ZN(n622) );
  XNOR2_X1 U723 ( .A(n666), .B(KEYINPUT105), .ZN(n731) );
  INV_X1 U724 ( .A(n731), .ZN(n679) );
  NOR2_X1 U725 ( .A1(n737), .A2(n679), .ZN(n623) );
  XNOR2_X1 U726 ( .A(n365), .B(G119), .ZN(G21) );
  XOR2_X1 U727 ( .A(KEYINPUT88), .B(KEYINPUT48), .Z(n656) );
  XOR2_X1 U728 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n629) );
  AND2_X1 U729 ( .A1(n630), .A2(n624), .ZN(n625) );
  NAND2_X1 U730 ( .A1(n630), .A2(n749), .ZN(n631) );
  INV_X1 U731 ( .A(KEYINPUT67), .ZN(n633) );
  INV_X1 U732 ( .A(n638), .ZN(n722) );
  INV_X1 U733 ( .A(n649), .ZN(n640) );
  NAND2_X1 U734 ( .A1(n640), .A2(n663), .ZN(n641) );
  NAND2_X1 U735 ( .A1(n644), .A2(n364), .ZN(n652) );
  NOR2_X1 U736 ( .A1(n646), .A2(n645), .ZN(n724) );
  INV_X1 U737 ( .A(n652), .ZN(n720) );
  INV_X1 U738 ( .A(n753), .ZN(n677) );
  NAND2_X1 U739 ( .A1(n720), .A2(n677), .ZN(n653) );
  NAND2_X1 U740 ( .A1(KEYINPUT47), .A2(n653), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n659), .A2(n724), .ZN(n660) );
  XOR2_X1 U742 ( .A(n660), .B(KEYINPUT110), .Z(n807) );
  INV_X1 U743 ( .A(n807), .ZN(n661) );
  INV_X1 U744 ( .A(KEYINPUT86), .ZN(n662) );
  INV_X1 U745 ( .A(n676), .ZN(n672) );
  INV_X1 U746 ( .A(n666), .ZN(n667) );
  AND2_X1 U747 ( .A1(n665), .A2(n667), .ZN(n668) );
  AND2_X1 U748 ( .A1(n737), .A2(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n716) );
  NAND2_X1 U750 ( .A1(n672), .A2(n745), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT31), .B(KEYINPUT101), .Z(n673) );
  XNOR2_X1 U752 ( .A(n674), .B(n673), .ZN(n725) );
  NAND2_X1 U753 ( .A1(n377), .A2(n665), .ZN(n675) );
  OR2_X1 U754 ( .A1(n725), .A2(n367), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U756 ( .A1(n737), .A2(n679), .ZN(n680) );
  OR2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n708) );
  NAND2_X1 U758 ( .A1(n683), .A2(n685), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n684), .A2(KEYINPUT85), .ZN(n689) );
  AND2_X1 U760 ( .A1(n685), .A2(KEYINPUT2), .ZN(n686) );
  NOR2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n688) );
  INV_X1 U762 ( .A(KEYINPUT2), .ZN(n730) );
  OR2_X1 U763 ( .A1(n807), .A2(n730), .ZN(n690) );
  XOR2_X1 U764 ( .A(KEYINPUT82), .B(n690), .Z(n691) );
  INV_X1 U765 ( .A(KEYINPUT78), .ZN(n692) );
  NAND2_X1 U766 ( .A1(n778), .A2(G472), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n694), .B(KEYINPUT62), .ZN(n695) );
  XNOR2_X1 U768 ( .A(n696), .B(n695), .ZN(n698) );
  INV_X1 U769 ( .A(G952), .ZN(n697) );
  NAND2_X1 U770 ( .A1(n698), .A2(n474), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n699), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U772 ( .A1(n778), .A2(G210), .ZN(n704) );
  XNOR2_X1 U773 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n700) );
  XOR2_X1 U774 ( .A(n700), .B(KEYINPUT55), .Z(n701) );
  XNOR2_X1 U775 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n705), .A2(n474), .ZN(n707) );
  XNOR2_X1 U777 ( .A(KEYINPUT87), .B(KEYINPUT56), .ZN(n706) );
  XNOR2_X1 U778 ( .A(n707), .B(n706), .ZN(G51) );
  XNOR2_X1 U779 ( .A(G101), .B(n708), .ZN(G3) );
  NAND2_X1 U780 ( .A1(n367), .A2(n722), .ZN(n709) );
  XNOR2_X1 U781 ( .A(n709), .B(G104), .ZN(G6) );
  XOR2_X1 U782 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n711) );
  XNOR2_X1 U783 ( .A(G107), .B(KEYINPUT26), .ZN(n710) );
  XNOR2_X1 U784 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(n712), .Z(n714) );
  NAND2_X1 U786 ( .A1(n367), .A2(n724), .ZN(n713) );
  XNOR2_X1 U787 ( .A(n714), .B(n713), .ZN(G9) );
  XOR2_X1 U788 ( .A(G110), .B(KEYINPUT113), .Z(n715) );
  XNOR2_X1 U789 ( .A(n716), .B(n715), .ZN(G12) );
  XOR2_X1 U790 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n718) );
  NAND2_X1 U791 ( .A1(n720), .A2(n724), .ZN(n717) );
  XNOR2_X1 U792 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U793 ( .A(G128), .B(n719), .ZN(G30) );
  NAND2_X1 U794 ( .A1(n720), .A2(n722), .ZN(n721) );
  XNOR2_X1 U795 ( .A(n721), .B(G146), .ZN(G48) );
  NAND2_X1 U796 ( .A1(n725), .A2(n722), .ZN(n723) );
  XNOR2_X1 U797 ( .A(n723), .B(G113), .ZN(G15) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U799 ( .A(n726), .B(G116), .ZN(G18) );
  XOR2_X1 U800 ( .A(G125), .B(KEYINPUT37), .Z(n727) );
  XNOR2_X1 U801 ( .A(n728), .B(n727), .ZN(G27) );
  NAND2_X1 U802 ( .A1(n732), .A2(n731), .ZN(n735) );
  XNOR2_X1 U803 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n733) );
  XNOR2_X1 U804 ( .A(n733), .B(KEYINPUT49), .ZN(n734) );
  XNOR2_X1 U805 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n736), .A2(n665), .ZN(n743) );
  XOR2_X1 U807 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n740) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U809 ( .A(n740), .B(n739), .ZN(n741) );
  XOR2_X1 U810 ( .A(KEYINPUT117), .B(n741), .Z(n742) );
  NOR2_X1 U811 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U812 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U813 ( .A(n746), .B(KEYINPUT51), .ZN(n748) );
  NAND2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n759) );
  NOR2_X1 U815 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U816 ( .A1(n752), .A2(n751), .ZN(n755) );
  NOR2_X1 U817 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U818 ( .A(KEYINPUT119), .B(n756), .ZN(n757) );
  NAND2_X1 U819 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U820 ( .A(KEYINPUT52), .B(n760), .Z(n761) );
  NOR2_X1 U821 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U822 ( .A(KEYINPUT121), .B(n764), .Z(n765) );
  NAND2_X1 U823 ( .A1(n387), .A2(G469), .ZN(n769) );
  XOR2_X1 U824 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n766) );
  NOR2_X1 U825 ( .A1(n781), .A2(n770), .ZN(G54) );
  NAND2_X1 U826 ( .A1(n778), .A2(G475), .ZN(n772) );
  XNOR2_X1 U827 ( .A(n772), .B(n534), .ZN(n773) );
  NAND2_X1 U828 ( .A1(n387), .A2(G478), .ZN(n776) );
  XNOR2_X1 U829 ( .A(n774), .B(KEYINPUT122), .ZN(n775) );
  XNOR2_X1 U830 ( .A(n776), .B(n775), .ZN(n777) );
  NOR2_X1 U831 ( .A1(n781), .A2(n777), .ZN(G63) );
  NAND2_X1 U832 ( .A1(n387), .A2(G217), .ZN(n780) );
  NAND2_X1 U833 ( .A1(G953), .A2(G224), .ZN(n782) );
  XNOR2_X1 U834 ( .A(KEYINPUT61), .B(n782), .ZN(n783) );
  NAND2_X1 U835 ( .A1(n783), .A2(G898), .ZN(n784) );
  NAND2_X1 U836 ( .A1(n785), .A2(n784), .ZN(n790) );
  XNOR2_X1 U837 ( .A(n363), .B(G101), .ZN(n788) );
  NOR2_X1 U838 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U839 ( .A(n790), .B(n789), .ZN(G69) );
  XOR2_X1 U840 ( .A(KEYINPUT125), .B(n791), .Z(n792) );
  XNOR2_X1 U841 ( .A(n793), .B(n792), .ZN(n794) );
  XOR2_X1 U842 ( .A(n795), .B(n794), .Z(n799) );
  XOR2_X1 U843 ( .A(n799), .B(n362), .Z(n798) );
  NAND2_X1 U844 ( .A1(n798), .A2(n797), .ZN(n804) );
  XNOR2_X1 U845 ( .A(n799), .B(G227), .ZN(n800) );
  XNOR2_X1 U846 ( .A(n800), .B(KEYINPUT126), .ZN(n801) );
  NAND2_X1 U847 ( .A1(n801), .A2(G900), .ZN(n802) );
  NAND2_X1 U848 ( .A1(G953), .A2(n802), .ZN(n803) );
  NAND2_X1 U849 ( .A1(n804), .A2(n803), .ZN(G72) );
  XNOR2_X1 U850 ( .A(G143), .B(n805), .ZN(G45) );
  XNOR2_X1 U851 ( .A(n361), .B(G131), .ZN(G33) );
  XOR2_X1 U852 ( .A(G134), .B(n807), .Z(G36) );
  XOR2_X1 U853 ( .A(n808), .B(G137), .Z(n809) );
  XNOR2_X1 U854 ( .A(KEYINPUT127), .B(n809), .ZN(G39) );
endmodule

