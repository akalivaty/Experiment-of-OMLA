

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  INV_X1 U325 ( .A(n525), .ZN(n516) );
  NOR2_X2 U326 ( .A1(n516), .A2(n471), .ZN(n559) );
  XNOR2_X1 U327 ( .A(n458), .B(n457), .ZN(n547) );
  XNOR2_X1 U328 ( .A(KEYINPUT48), .B(n466), .ZN(n540) );
  AND2_X1 U329 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U330 ( .A(n358), .B(n357), .ZN(n361) );
  XNOR2_X1 U331 ( .A(KEYINPUT38), .B(n449), .ZN(n496) );
  XOR2_X1 U332 ( .A(n469), .B(KEYINPUT28), .Z(n521) );
  XNOR2_X1 U333 ( .A(n396), .B(n364), .ZN(n514) );
  OR2_X1 U334 ( .A1(n371), .A2(n564), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n402), .B(n422), .ZN(n403) );
  INV_X1 U336 ( .A(KEYINPUT94), .ZN(n355) );
  XNOR2_X1 U337 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U338 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U339 ( .A(n389), .B(n388), .ZN(n390) );
  OR2_X1 U340 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U341 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U342 ( .A(n374), .B(KEYINPUT97), .ZN(n478) );
  XNOR2_X1 U343 ( .A(n409), .B(n408), .ZN(n577) );
  INV_X1 U344 ( .A(G36GAT), .ZN(n450) );
  XNOR2_X1 U345 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U346 ( .A(n450), .B(KEYINPUT104), .ZN(n451) );
  XNOR2_X1 U347 ( .A(n475), .B(n474), .ZN(G1349GAT) );
  XNOR2_X1 U348 ( .A(n452), .B(n451), .ZN(G1329GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n412) );
  XOR2_X1 U350 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n295) );
  XNOR2_X1 U351 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n313) );
  XOR2_X1 U353 ( .A(G155GAT), .B(G162GAT), .Z(n297) );
  XNOR2_X1 U354 ( .A(G127GAT), .B(G148GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U356 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n299) );
  XNOR2_X1 U357 ( .A(G1GAT), .B(G57GAT), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U359 ( .A(n301), .B(n300), .Z(n311) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n302), .B(G120GAT), .ZN(n341) );
  XOR2_X1 U362 ( .A(KEYINPUT5), .B(n341), .Z(n304) );
  NAND2_X1 U363 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U365 ( .A(G134GAT), .B(KEYINPUT78), .Z(n381) );
  XOR2_X1 U366 ( .A(G85GAT), .B(n381), .Z(n307) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n305) );
  XNOR2_X1 U368 ( .A(n305), .B(KEYINPUT2), .ZN(n327) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(n327), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n563) );
  XOR2_X1 U374 ( .A(KEYINPUT88), .B(G218GAT), .Z(n315) );
  XOR2_X1 U375 ( .A(G197GAT), .B(KEYINPUT21), .Z(n359) );
  XOR2_X1 U376 ( .A(G22GAT), .B(G155GAT), .Z(n399) );
  XNOR2_X1 U377 ( .A(n359), .B(n399), .ZN(n314) );
  XNOR2_X1 U378 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .Z(n388) );
  XOR2_X1 U380 ( .A(n316), .B(n388), .Z(n321) );
  XOR2_X1 U381 ( .A(KEYINPUT22), .B(G204GAT), .Z(n318) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U384 ( .A(KEYINPUT24), .B(n319), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U386 ( .A(KEYINPUT89), .B(G211GAT), .Z(n323) );
  XNOR2_X1 U387 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U389 ( .A(n325), .B(n324), .Z(n329) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n326), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U392 ( .A(n415), .B(n327), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n469) );
  XOR2_X1 U394 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n331) );
  XNOR2_X1 U395 ( .A(G190GAT), .B(G134GAT), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U397 ( .A(n332), .B(G99GAT), .Z(n334) );
  XOR2_X1 U398 ( .A(G15GAT), .B(G127GAT), .Z(n400) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(n400), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U401 ( .A(G183GAT), .B(KEYINPUT86), .Z(n336) );
  XNOR2_X1 U402 ( .A(G71GAT), .B(KEYINPUT85), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U404 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U405 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n340) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n340), .B(n339), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n341), .B(n352), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U410 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n345) );
  NAND2_X1 U411 ( .A1(G227GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U412 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U413 ( .A(G176GAT), .B(n346), .Z(n347) );
  XOR2_X1 U414 ( .A(n348), .B(n347), .Z(n525) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G183GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n349), .B(G211GAT), .ZN(n396) );
  XOR2_X1 U417 ( .A(G64GAT), .B(G92GAT), .Z(n351) );
  XNOR2_X1 U418 ( .A(G176GAT), .B(G204GAT), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n423) );
  XNOR2_X1 U420 ( .A(n352), .B(n423), .ZN(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT79), .B(G218GAT), .Z(n354) );
  XNOR2_X1 U422 ( .A(G36GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n382) );
  XOR2_X1 U424 ( .A(n382), .B(KEYINPUT95), .Z(n358) );
  NAND2_X1 U425 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n359), .B(KEYINPUT93), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  NOR2_X1 U429 ( .A1(n516), .A2(n514), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n365), .B(KEYINPUT96), .ZN(n366) );
  NOR2_X1 U431 ( .A1(n469), .A2(n366), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n367), .B(KEYINPUT25), .ZN(n369) );
  XNOR2_X1 U433 ( .A(KEYINPUT27), .B(n514), .ZN(n371) );
  NAND2_X1 U434 ( .A1(n516), .A2(n469), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n368), .B(KEYINPUT26), .ZN(n564) );
  AND2_X1 U436 ( .A1(n369), .A2(n293), .ZN(n370) );
  NOR2_X1 U437 ( .A1(n563), .A2(n370), .ZN(n373) );
  INV_X1 U438 ( .A(n563), .ZN(n512) );
  NOR2_X1 U439 ( .A1(n512), .A2(n371), .ZN(n542) );
  NAND2_X1 U440 ( .A1(n542), .A2(n521), .ZN(n524) );
  NOR2_X1 U441 ( .A1(n525), .A2(n524), .ZN(n372) );
  XOR2_X1 U442 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n376) );
  XNOR2_X1 U443 ( .A(G43GAT), .B(G29GAT), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U445 ( .A(KEYINPUT69), .B(n377), .Z(n435) );
  XOR2_X1 U446 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n379) );
  XNOR2_X1 U447 ( .A(G106GAT), .B(G92GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n435), .B(n380), .ZN(n393) );
  XOR2_X1 U450 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U451 ( .A1(G232GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n391) );
  XOR2_X1 U453 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n386) );
  XNOR2_X1 U454 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U456 ( .A(G99GAT), .B(G85GAT), .Z(n413) );
  XOR2_X1 U457 ( .A(n387), .B(n413), .Z(n389) );
  XOR2_X1 U458 ( .A(n393), .B(n392), .Z(n560) );
  XOR2_X1 U459 ( .A(n560), .B(KEYINPUT36), .Z(n583) );
  NOR2_X1 U460 ( .A1(n478), .A2(n583), .ZN(n410) );
  XOR2_X1 U461 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n395) );
  XNOR2_X1 U462 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n396), .B(KEYINPUT14), .ZN(n398) );
  AND2_X1 U465 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n404) );
  XOR2_X1 U467 ( .A(n400), .B(n399), .Z(n402) );
  XNOR2_X1 U468 ( .A(G71GAT), .B(G57GAT), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n401), .B(KEYINPUT13), .ZN(n422) );
  XNOR2_X1 U470 ( .A(n405), .B(G64GAT), .ZN(n407) );
  XOR2_X1 U471 ( .A(KEYINPUT70), .B(G1GAT), .Z(n431) );
  XOR2_X1 U472 ( .A(n431), .B(G78GAT), .Z(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  NAND2_X1 U474 ( .A1(n410), .A2(n577), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n511) );
  XNOR2_X1 U476 ( .A(G120GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n414), .B(KEYINPUT75), .ZN(n427) );
  XOR2_X1 U478 ( .A(n415), .B(KEYINPUT31), .Z(n417) );
  NAND2_X1 U479 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U481 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n419) );
  XNOR2_X1 U482 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U484 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n457) );
  INV_X1 U488 ( .A(n457), .ZN(n573) );
  XOR2_X1 U489 ( .A(G113GAT), .B(G15GAT), .Z(n429) );
  XNOR2_X1 U490 ( .A(G36GAT), .B(G50GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U492 ( .A(n430), .B(G197GAT), .Z(n433) );
  XNOR2_X1 U493 ( .A(G169GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n448) );
  XOR2_X1 U496 ( .A(KEYINPUT65), .B(G8GAT), .Z(n437) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(G141GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U499 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n439) );
  XNOR2_X1 U500 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U503 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n443) );
  NAND2_X1 U504 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U506 ( .A(KEYINPUT71), .B(n444), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U508 ( .A(n448), .B(n447), .Z(n543) );
  NOR2_X1 U509 ( .A1(n573), .A2(n543), .ZN(n479) );
  NAND2_X1 U510 ( .A1(n511), .A2(n479), .ZN(n449) );
  NOR2_X1 U511 ( .A1(n496), .A2(n514), .ZN(n452) );
  INV_X1 U512 ( .A(n543), .ZN(n568) );
  NOR2_X1 U513 ( .A1(n577), .A2(n583), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT45), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n454), .A2(n457), .ZN(n455) );
  NOR2_X1 U516 ( .A1(n568), .A2(n455), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT113), .ZN(n465) );
  XNOR2_X1 U518 ( .A(KEYINPUT111), .B(n577), .ZN(n557) );
  INV_X1 U519 ( .A(KEYINPUT41), .ZN(n458) );
  NOR2_X1 U520 ( .A1(n543), .A2(n547), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n459), .B(KEYINPUT46), .ZN(n460) );
  NOR2_X1 U522 ( .A1(n557), .A2(n460), .ZN(n461) );
  XOR2_X1 U523 ( .A(KEYINPUT112), .B(n461), .Z(n462) );
  NOR2_X1 U524 ( .A1(n560), .A2(n462), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n463), .B(KEYINPUT47), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n540), .A2(n514), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT54), .ZN(n566) );
  NAND2_X1 U528 ( .A1(n566), .A2(n512), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT55), .ZN(n471) );
  INV_X1 U531 ( .A(n547), .ZN(n529) );
  NAND2_X1 U532 ( .A1(n559), .A2(n529), .ZN(n475) );
  XOR2_X1 U533 ( .A(G176GAT), .B(KEYINPUT57), .Z(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n472) );
  NOR2_X1 U535 ( .A1(n560), .A2(n577), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(n476), .Z(n477) );
  NOR2_X1 U537 ( .A1(n478), .A2(n477), .ZN(n499) );
  NAND2_X1 U538 ( .A1(n479), .A2(n499), .ZN(n488) );
  NOR2_X1 U539 ( .A1(n512), .A2(n488), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n482), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n514), .A2(n488), .ZN(n484) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  NOR2_X1 U546 ( .A1(n516), .A2(n488), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n521), .A2(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(G1327GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n492) );
  NOR2_X1 U554 ( .A1(n512), .A2(n496), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n496), .A2(n516), .ZN(n494) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n521), .A2(n496), .ZN(n497) );
  XOR2_X1 U561 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  NAND2_X1 U562 ( .A1(n543), .A2(n529), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(KEYINPUT105), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n510), .A2(n499), .ZN(n507) );
  NOR2_X1 U565 ( .A1(n512), .A2(n507), .ZN(n501) );
  XNOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n507), .ZN(n503) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n516), .A2(n507), .ZN(n505) );
  XNOR2_X1 U572 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n521), .A2(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n512), .A2(n520), .ZN(n513) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n520), .ZN(n517) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(n523), .B(n522), .Z(G1339GAT) );
  NOR2_X1 U590 ( .A1(n540), .A2(n524), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT114), .B(n527), .Z(n536) );
  NAND2_X1 U593 ( .A1(n536), .A2(n568), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U596 ( .A1(n529), .A2(n536), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U600 ( .A1(n557), .A2(n536), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U602 ( .A(G127GAT), .B(n535), .Z(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U604 ( .A1(n536), .A2(n560), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  NOR2_X1 U607 ( .A1(n564), .A2(n540), .ZN(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n553) );
  NOR2_X1 U609 ( .A1(n543), .A2(n553), .ZN(n544) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n547), .A2(n553), .ZN(n548) );
  XOR2_X1 U615 ( .A(n549), .B(n548), .Z(G1345GAT) );
  NOR2_X1 U616 ( .A1(n577), .A2(n553), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  INV_X1 U620 ( .A(n560), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n568), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n557), .A2(n559), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT58), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n562), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  AND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT122), .B(n567), .Z(n584) );
  INV_X1 U634 ( .A(n584), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n568), .A2(n572), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n579) );
  OR2_X1 U643 ( .A1(n577), .A2(n584), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

