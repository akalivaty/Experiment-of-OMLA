//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT64), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G226), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G97), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n256), .A2(new_n258), .A3(new_n262), .A4(new_n259), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n250), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n261), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(G274), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n265), .A2(new_n269), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT66), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n272), .B2(G238), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n267), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G169), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT14), .ZN(new_n280));
  INV_X1    g0080(.A(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G179), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n278), .A2(new_n283), .A3(G169), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n215), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n250), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n225), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n292), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n287), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT11), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT12), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n302), .B2(new_n219), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n304));
  INV_X1    g0104(.A(new_n287), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G1), .B2(new_n207), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n303), .A2(new_n304), .B1(new_n219), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n294), .A2(new_n295), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n297), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n285), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n281), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n278), .A2(KEYINPUT72), .A3(G200), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n309), .B1(new_n278), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n270), .B1(new_n272), .B2(G226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n257), .A2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n324), .B1(new_n225), .B2(new_n257), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(G222), .B2(new_n255), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n322), .B1(new_n265), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n301), .A2(new_n202), .ZN(new_n329));
  INV_X1    g0129(.A(new_n306), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n202), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT68), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n291), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT67), .ZN(new_n334));
  INV_X1    g0134(.A(G58), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT8), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n338), .B2(KEYINPUT67), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n333), .B1(new_n339), .B2(new_n289), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n287), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n327), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n328), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT9), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n343), .B(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT10), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n327), .A2(new_n317), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(G200), .B2(new_n327), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n349), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n339), .A2(new_n301), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n330), .B2(new_n339), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT78), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT75), .B1(new_n335), .B2(new_n219), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT75), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(G58), .A3(G68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n201), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n291), .A2(G159), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G20), .B1(new_n251), .B2(new_n253), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT76), .B1(new_n367), .B2(KEYINPUT7), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT76), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n370), .C1(new_n257), .C2(G20), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n253), .B1(new_n372), .B2(G33), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n370), .A2(G20), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n368), .A2(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n366), .B1(new_n375), .B2(new_n219), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT77), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n252), .A2(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n384), .A3(G33), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(KEYINPUT3), .B2(new_n250), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n382), .A2(new_n384), .A3(new_n386), .A4(G33), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n207), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT7), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n390), .B2(KEYINPUT7), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT16), .B(new_n366), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n394), .A2(new_n287), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n359), .B1(new_n381), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n324), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G226), .B2(new_n397), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n388), .B2(new_n389), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n250), .A2(new_n221), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n266), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n270), .B1(G232), .B2(new_n271), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n404), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n407), .A2(G169), .B1(G179), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT18), .B1(new_n396), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n364), .A2(new_n365), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n373), .A2(new_n374), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n254), .A2(new_n207), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n369), .B1(new_n413), .B2(new_n370), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n367), .A2(KEYINPUT76), .A3(KEYINPUT7), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(G68), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT77), .B1(new_n417), .B2(KEYINPUT16), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n287), .A3(new_n394), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n358), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n408), .A2(G179), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n405), .A2(new_n406), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n345), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n313), .B1(new_n405), .B2(new_n406), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n402), .A2(new_n317), .A3(new_n404), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n420), .A3(new_n358), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n429), .A2(new_n420), .A3(KEYINPUT17), .A4(new_n358), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n410), .A2(new_n426), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n270), .B1(new_n272), .B2(G244), .ZN(new_n435));
  OR2_X1    g0235(.A1(KEYINPUT69), .A2(G107), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT69), .A2(G107), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n323), .A2(new_n220), .B1(new_n438), .B2(new_n257), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(G232), .B2(new_n255), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n435), .B1(new_n265), .B2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(G179), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n302), .A2(new_n225), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n306), .B2(new_n225), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n338), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT70), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(new_n289), .ZN(new_n448));
  INV_X1    g0248(.A(new_n447), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT70), .A3(new_n288), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n445), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n444), .B1(new_n287), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n441), .B2(new_n345), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n441), .A2(G200), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n452), .C1(new_n317), .C2(new_n441), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n321), .A2(new_n355), .A3(new_n434), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n286), .A2(new_n215), .B1(G20), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n207), .C1(G33), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(KEYINPUT20), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n461), .B2(new_n464), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n301), .A2(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n206), .A2(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n305), .A2(new_n301), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(G116), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n466), .A2(new_n467), .ZN(new_n476));
  INV_X1    g0276(.A(new_n469), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n471), .B2(new_n460), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT85), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n481), .A2(new_n265), .A3(G274), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(new_n265), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n489), .B2(G270), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n388), .A2(new_n389), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G257), .A2(G1698), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n228), .B2(G1698), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(new_n493), .B1(G303), .B2(new_n254), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n490), .B1(new_n494), .B2(new_n265), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n480), .A2(G169), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n480), .A2(KEYINPUT21), .A3(new_n495), .A4(G169), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n490), .B(G179), .C1(new_n494), .C2(new_n265), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n480), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n480), .B1(G200), .B2(new_n495), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n317), .B2(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G238), .A2(G1698), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n226), .B2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n251), .A2(KEYINPUT74), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(G33), .B2(new_n372), .ZN(new_n511));
  INV_X1    g0311(.A(new_n389), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n265), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n483), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT83), .B1(new_n268), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT83), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n265), .A2(new_n518), .A3(G274), .A4(new_n483), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n266), .A2(new_n222), .A3(new_n483), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G200), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n302), .A2(new_n447), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n491), .A2(new_n207), .A3(G68), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n259), .B2(new_n207), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n436), .A2(new_n463), .A3(new_n437), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT84), .B(G87), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n528), .B1(new_n289), .B2(new_n463), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n526), .B1(new_n535), .B2(new_n287), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n472), .A2(G87), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n521), .B1(new_n517), .B2(new_n519), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n491), .A2(new_n509), .B1(G33), .B2(G116), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(G190), .C1(new_n539), .C2(new_n265), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n524), .A2(new_n536), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n472), .A2(new_n449), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n532), .A2(new_n533), .ZN(new_n543));
  AOI21_X1  g0343(.A(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(G68), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n525), .B(new_n542), .C1(new_n545), .C2(new_n305), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n345), .B1(new_n515), .B2(new_n523), .ZN(new_n547));
  INV_X1    g0347(.A(G179), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n538), .B(new_n548), .C1(new_n539), .C2(new_n265), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n507), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n227), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  XOR2_X1   g0353(.A(G97), .B(G107), .Z(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(KEYINPUT6), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n375), .B2(new_n438), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n287), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n302), .A2(new_n463), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n471), .B2(new_n463), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n488), .A2(G257), .A3(new_n265), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT80), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(new_n484), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n563), .B2(new_n484), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n397), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n462), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n226), .A2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n511), .B2(new_n512), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n567), .B1(new_n574), .B2(new_n265), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n345), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n567), .B(new_n548), .C1(new_n574), .C2(new_n265), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n562), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT82), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n567), .B(KEYINPUT81), .C1(new_n574), .C2(new_n265), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(G200), .A4(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n567), .B(G190), .C1(new_n574), .C2(new_n265), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n584), .A2(new_n558), .A3(new_n561), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n313), .B1(new_n575), .B2(new_n579), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n581), .B1(new_n587), .B2(new_n582), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n578), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n489), .A2(G264), .ZN(new_n590));
  MUX2_X1   g0390(.A(G250), .B(G257), .S(G1698), .Z(new_n591));
  AOI22_X1  g0391(.A1(new_n491), .A2(new_n591), .B1(G33), .B2(G294), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n484), .B(new_n590), .C1(new_n592), .C2(new_n265), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n313), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT88), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n596), .A3(new_n313), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n593), .A2(G190), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g0399(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n600));
  NOR4_X1   g0400(.A1(new_n600), .A2(new_n254), .A3(G20), .A4(new_n221), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n207), .B(G87), .C1(new_n511), .C2(new_n512), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(KEYINPUT22), .ZN(new_n603));
  OR3_X1    g0403(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n289), .B2(new_n460), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n438), .A2(G20), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(KEYINPUT23), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT87), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT22), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n544), .B2(G87), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n607), .C1(new_n612), .C2(new_n601), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(KEYINPUT24), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT87), .B(new_n615), .C1(new_n603), .C2(new_n608), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n287), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n300), .A2(G20), .A3(new_n227), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT25), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(G107), .B2(new_n472), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n599), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n589), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n609), .A2(KEYINPUT24), .A3(new_n613), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(new_n287), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n593), .A2(new_n345), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G179), .B2(new_n593), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n552), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n459), .A2(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n347), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n318), .B1(new_n314), .B2(new_n315), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n311), .B1(new_n633), .B2(new_n454), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n432), .A3(new_n433), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n410), .A2(new_n426), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT93), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n353), .A2(new_n354), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n638), .B2(KEYINPUT93), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n632), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT91), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n578), .B(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n541), .A2(new_n550), .A3(KEYINPUT89), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT89), .B1(new_n541), .B2(new_n550), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT26), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n551), .A2(new_n578), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT26), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n558), .A2(new_n561), .B1(new_n575), .B2(new_n345), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(new_n577), .A3(new_n550), .A4(new_n541), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT92), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n550), .B1(new_n649), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n627), .B1(new_n617), .B2(new_n620), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n648), .B1(new_n660), .B2(new_n503), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n580), .A2(G200), .A3(new_n582), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT82), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n583), .A3(new_n585), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n599), .A2(new_n617), .A3(new_n620), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n578), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n659), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n551), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n541), .A2(new_n550), .A3(KEYINPUT89), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n629), .B2(new_n504), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n622), .A3(KEYINPUT90), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n658), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n643), .B1(new_n459), .B2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n300), .A2(new_n207), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n480), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT94), .Z(new_n683));
  OR2_X1    g0483(.A1(new_n507), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n503), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n681), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n617), .B2(new_n620), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n629), .B1(new_n621), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n660), .A2(new_n691), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n504), .A2(new_n681), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n694), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n210), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n530), .A2(new_n531), .A3(G116), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n213), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n515), .A2(new_n523), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n575), .A3(new_n593), .A4(new_n495), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n575), .A2(new_n500), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n592), .A2(new_n265), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n714), .A3(new_n590), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT95), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n712), .B1(new_n719), .B2(KEYINPUT30), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  AOI211_X1 g0521(.A(new_n721), .B(new_n713), .C1(new_n717), .C2(new_n718), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n681), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT31), .B(new_n681), .C1(new_n720), .C2(new_n722), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n725), .B(new_n726), .C1(new_n630), .C2(new_n681), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n673), .A2(new_n667), .ZN(new_n730));
  INV_X1    g0530(.A(new_n550), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n645), .A2(new_n648), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n655), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n652), .A2(new_n656), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n681), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT96), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT96), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n738), .B(new_n739), .C1(new_n674), .C2(new_n681), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n732), .A2(KEYINPUT26), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n731), .B1(new_n650), .B2(new_n655), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n742), .B(new_n743), .C1(new_n666), .C2(new_n661), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n729), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n709), .B1(new_n746), .B2(G1), .ZN(G364));
  NOR2_X1   g0547(.A1(new_n299), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n206), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n704), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n687), .A2(new_n688), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n690), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n703), .A2(new_n254), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G355), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G116), .B2(new_n210), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n244), .A2(G45), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n491), .A2(new_n703), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n482), .B2(new_n214), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n215), .B1(G20), .B2(new_n345), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n751), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G329), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(new_n548), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n776), .A2(new_n313), .A3(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT33), .B(G317), .Z(new_n779));
  OAI21_X1  g0579(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n776), .A2(new_n317), .A3(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n257), .B1(new_n781), .B2(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n775), .A2(new_n771), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n780), .B(new_n785), .C1(G311), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n776), .A2(new_n317), .A3(new_n313), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G326), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n317), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n207), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n770), .A2(new_n317), .A3(G200), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT97), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT97), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n795), .A2(KEYINPUT98), .B1(new_n800), .B2(G283), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n788), .B(new_n801), .C1(KEYINPUT98), .C2(new_n795), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n778), .A2(new_n219), .B1(new_n786), .B2(new_n225), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G50), .B2(new_n789), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(G107), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n772), .A2(KEYINPUT32), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n794), .A2(new_n463), .ZN(new_n808));
  INV_X1    g0608(.A(new_n784), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n808), .C1(new_n531), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT32), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n773), .B2(G159), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n254), .B(new_n812), .C1(G58), .C2(new_n781), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n804), .A2(new_n805), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n802), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n769), .B1(new_n815), .B2(new_n766), .ZN(new_n816));
  INV_X1    g0616(.A(new_n765), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n686), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n754), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT99), .ZN(G396));
  OAI21_X1  g0620(.A(new_n456), .B1(new_n452), .B2(new_n691), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n454), .ZN(new_n822));
  INV_X1    g0622(.A(new_n454), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n691), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n736), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n751), .B1(new_n827), .B2(new_n728), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n728), .B2(new_n827), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  INV_X1    g0630(.A(new_n781), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n778), .B1(new_n831), .B2(new_n792), .ZN(new_n832));
  INV_X1    g0632(.A(G311), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n790), .A2(new_n783), .B1(new_n772), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n800), .A2(G87), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n809), .A2(G107), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n257), .B(new_n808), .C1(G116), .C2(new_n787), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n777), .A2(G150), .B1(G159), .B2(new_n787), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT100), .B(G143), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n841), .B2(new_n790), .C1(new_n831), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n843), .A2(new_n844), .B1(G68), .B2(new_n800), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n809), .A2(G50), .B1(new_n773), .B2(G132), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(new_n491), .C1(new_n335), .C2(new_n794), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n766), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n766), .A2(new_n763), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n752), .B1(new_n225), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(new_n826), .C2(new_n764), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n829), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  OR2_X1    g0655(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n856), .A2(G116), .A3(new_n216), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT36), .Z(new_n859));
  NAND4_X1  g0659(.A1(new_n214), .A2(new_n360), .A3(G77), .A4(new_n362), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n202), .A2(G68), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n206), .B(G13), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n748), .A2(new_n206), .ZN(new_n864));
  INV_X1    g0664(.A(new_n824), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n736), .B2(new_n826), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n309), .A2(new_n691), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n311), .A2(new_n320), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n310), .B(new_n681), .C1(new_n633), .C2(new_n285), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n679), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n392), .A2(new_n393), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n378), .B1(new_n875), .B2(new_n411), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n359), .B1(new_n395), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n434), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n409), .B2(new_n679), .ZN(new_n880));
  INV_X1    g0680(.A(new_n430), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n421), .A2(new_n424), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n421), .A2(new_n874), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n430), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n879), .A2(new_n887), .A3(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n873), .A2(new_n892), .B1(new_n636), .B2(new_n679), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n285), .A2(new_n310), .A3(new_n691), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n891), .ZN(new_n896));
  INV_X1    g0696(.A(new_n891), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n434), .A2(new_n421), .A3(new_n874), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT102), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT102), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n434), .A2(new_n900), .A3(new_n421), .A4(new_n874), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n883), .A2(new_n884), .A3(new_n430), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(KEYINPUT101), .A3(new_n886), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT101), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n899), .A2(new_n901), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n897), .B1(new_n907), .B2(new_n889), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n895), .B(new_n896), .C1(new_n908), .C2(KEYINPUT39), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n458), .A2(new_n745), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n737), .B2(new_n740), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT103), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(KEYINPUT103), .B(new_n911), .C1(new_n737), .C2(new_n740), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n643), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n910), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT104), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n825), .B1(new_n869), .B2(new_n870), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n727), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT40), .B1(new_n908), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n727), .A2(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(KEYINPUT40), .C2(new_n892), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n458), .A2(new_n727), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n927), .A2(new_n928), .A3(new_n688), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n864), .B1(new_n917), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n930), .A2(new_n931), .B1(new_n917), .B2(new_n929), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n863), .B1(new_n932), .B2(new_n933), .ZN(G367));
  OAI221_X1 g0734(.A(new_n767), .B1(new_n210), .B2(new_n447), .C1(new_n760), .C2(new_n239), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(new_n751), .ZN(new_n936));
  INV_X1    g0736(.A(new_n766), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n254), .B1(new_n800), .B2(G77), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT110), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n787), .A2(G50), .ZN(new_n940));
  AOI22_X1  g0740(.A1(G150), .A2(new_n781), .B1(new_n777), .B2(G159), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n790), .A2(new_n842), .B1(new_n772), .B2(new_n841), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n794), .A2(new_n219), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n784), .A2(new_n335), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n938), .A2(KEYINPUT110), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n794), .A2(new_n438), .B1(new_n786), .B2(new_n830), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT109), .Z(new_n949));
  AOI22_X1  g0749(.A1(G294), .A2(new_n777), .B1(new_n781), .B2(G303), .ZN(new_n950));
  INV_X1    g0750(.A(new_n491), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n789), .A2(G311), .B1(G317), .B2(new_n773), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n800), .A2(G97), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n809), .A2(G116), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT46), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n946), .A2(new_n947), .B1(new_n949), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n536), .A2(new_n537), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n681), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n550), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n648), .B2(new_n962), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n936), .B1(new_n937), .B2(new_n960), .C1(new_n965), .C2(new_n817), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n562), .A2(new_n681), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n664), .A2(new_n578), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n653), .A2(new_n577), .A3(new_n681), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n971), .A2(new_n695), .A3(new_n699), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n578), .B1(new_n968), .B2(new_n629), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n691), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n964), .B1(new_n978), .B2(KEYINPUT106), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n977), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT106), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n981), .A3(new_n965), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n979), .A2(KEYINPUT43), .A3(new_n980), .A4(new_n982), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n697), .A2(new_n971), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n701), .A2(new_n970), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  XOR2_X1   g0792(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n701), .B2(new_n970), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n700), .A2(new_n971), .A3(new_n993), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n696), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(KEYINPUT108), .B(new_n696), .C1(new_n992), .C2(new_n997), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n992), .A2(new_n696), .A3(new_n997), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n695), .B(new_n698), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n689), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n746), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n704), .B(KEYINPUT41), .Z(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n750), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n966), .B1(new_n990), .B2(new_n1009), .ZN(G387));
  INV_X1    g0810(.A(new_n1005), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n705), .B1(new_n746), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n746), .B2(new_n1011), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n236), .A2(new_n482), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1014), .A2(new_n759), .B1(new_n707), .B2(new_n755), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n337), .A2(G50), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT50), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n482), .B1(new_n219), .B2(new_n225), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n707), .B(new_n1018), .C1(new_n1017), .C2(new_n1016), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1015), .A2(new_n1019), .B1(G107), .B2(new_n210), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n752), .B1(new_n1020), .B2(new_n767), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n789), .A2(G159), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT112), .Z(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n491), .C1(new_n339), .C2(new_n778), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n831), .A2(new_n202), .B1(new_n786), .B2(new_n219), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G150), .B2(new_n773), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n794), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1028), .A2(new_n449), .B1(new_n809), .B2(G77), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1025), .A2(new_n954), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT113), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n1028), .A2(G283), .B1(new_n809), .B2(G294), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT114), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n781), .A2(G317), .B1(new_n789), .B2(G322), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n777), .A2(G311), .B1(G303), .B2(new_n787), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1035), .B1(new_n1038), .B2(KEYINPUT48), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1034), .B(new_n1039), .C1(KEYINPUT48), .C2(new_n1038), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n951), .B1(new_n791), .B2(new_n772), .C1(new_n799), .C2(new_n460), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n1040), .B2(KEYINPUT49), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1031), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1021), .B1(new_n1044), .B2(new_n937), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n695), .B2(new_n765), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1011), .B2(new_n750), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1013), .A2(new_n1047), .ZN(G393));
  NAND3_X1  g0848(.A1(new_n1002), .A2(new_n750), .A3(new_n998), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n248), .A2(new_n760), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n767), .B1(new_n463), .B2(new_n210), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n751), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n781), .A2(G159), .B1(new_n789), .B2(G150), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n836), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n794), .A2(new_n225), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G68), .B2(new_n809), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n777), .A2(G50), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n842), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n338), .A2(new_n787), .B1(new_n773), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n491), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n781), .A2(G311), .B1(new_n789), .B2(G317), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT52), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n257), .B1(new_n787), .B2(G294), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n777), .A2(G303), .B1(G322), .B2(new_n773), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1028), .A2(G116), .B1(new_n809), .B2(G283), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n805), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1055), .A2(new_n1061), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1052), .B1(new_n1068), .B2(new_n766), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n970), .B2(new_n817), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1049), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n746), .A2(new_n1011), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1003), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1073), .A2(new_n705), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1002), .A2(new_n998), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1072), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1071), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(G390));
  OAI22_X1  g0878(.A1(new_n778), .A2(new_n438), .B1(new_n790), .B2(new_n830), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n831), .A2(new_n460), .B1(new_n772), .B2(new_n792), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n254), .B1(new_n786), .B2(new_n463), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1082), .B(new_n1056), .C1(G87), .C2(new_n809), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G68), .B2(new_n800), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n781), .A2(G132), .B1(new_n789), .B2(G128), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n777), .A2(G137), .B1(G125), .B2(new_n773), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(G150), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n784), .A2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT53), .Z(new_n1091));
  NOR2_X1   g0891(.A1(new_n799), .A2(new_n202), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n257), .B1(new_n786), .B2(new_n1093), .C1(new_n794), .C2(new_n806), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n766), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n752), .B1(new_n339), .B2(new_n851), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n896), .B1(new_n908), .B2(KEYINPUT39), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n763), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n894), .B1(new_n866), .B2(new_n872), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n907), .A2(new_n889), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n891), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n744), .A2(new_n691), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n865), .B1(new_n1105), .B2(new_n822), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n894), .C1(new_n872), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n727), .A2(G330), .A3(new_n826), .A4(new_n871), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1102), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1100), .B1(new_n1114), .B2(new_n750), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n729), .A2(new_n458), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n643), .B(new_n1116), .C1(new_n914), .C2(new_n915), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n872), .B1(new_n728), .B2(new_n825), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n866), .B1(new_n1118), .B2(new_n1109), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT115), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n826), .B1(new_n728), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT115), .B1(new_n727), .B2(G330), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n872), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n704), .B1(new_n1114), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1115), .B1(new_n1127), .B2(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(KEYINPUT120), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1117), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1113), .B2(new_n1125), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n925), .A2(G330), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1135));
  NOR2_X1   g0935(.A1(new_n355), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n344), .A2(new_n874), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT119), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n355), .A2(new_n1135), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n925), .A2(new_n1145), .A3(G330), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n910), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n893), .A2(new_n909), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1145), .B1(new_n925), .B2(G330), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n688), .B(new_n1143), .C1(new_n921), .C2(new_n924), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1133), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1131), .B1(new_n1153), .B2(KEYINPUT57), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1133), .A2(KEYINPUT57), .A3(new_n1152), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1155), .A2(new_n704), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT57), .B1(new_n1133), .B2(new_n1152), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1143), .A2(new_n763), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n777), .A2(G132), .B1(new_n789), .B2(G125), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n781), .A2(G128), .B1(G137), .B2(new_n787), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n1089), .B2(new_n794), .C1(new_n784), .C2(new_n1093), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n773), .C2(G124), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n799), .B2(new_n806), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1164), .B2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n951), .A2(new_n264), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G50), .B1(new_n250), .B2(new_n264), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1165), .A2(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n943), .B1(G116), .B2(new_n789), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT117), .Z(new_n1173));
  AOI22_X1  g0973(.A1(new_n777), .A2(G97), .B1(new_n449), .B2(new_n787), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT116), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n831), .A2(new_n227), .B1(new_n772), .B2(new_n830), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G77), .B2(new_n809), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n799), .A2(new_n335), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n1169), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1173), .A2(new_n1175), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1171), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n766), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n752), .B(new_n1186), .C1(new_n202), .C2(new_n851), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1152), .A2(new_n750), .B1(new_n1160), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1159), .A2(new_n1188), .ZN(G375));
  INV_X1    g0989(.A(new_n1126), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1008), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n752), .B1(new_n219), .B2(new_n851), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n254), .B1(new_n438), .B2(new_n786), .C1(new_n447), .C2(new_n794), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n778), .A2(new_n460), .B1(new_n790), .B2(new_n792), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(G283), .C2(new_n781), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n784), .A2(new_n463), .B1(new_n772), .B2(new_n783), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT121), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(new_n225), .C2(new_n799), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n789), .A2(G132), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1089), .B2(new_n786), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n951), .B(new_n1201), .C1(G128), .C2(new_n773), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n841), .A2(new_n831), .B1(new_n778), .B2(new_n1093), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G50), .B2(new_n1028), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n806), .C2(new_n784), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1199), .B1(new_n1205), .B2(new_n1178), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT122), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n766), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1193), .B1(new_n1207), .B2(new_n1209), .C1(new_n871), .C2(new_n764), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1125), .B2(new_n749), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1192), .A2(new_n1212), .ZN(G381));
  INV_X1    g1013(.A(G378), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1159), .A2(new_n1214), .A3(new_n1188), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1077), .A2(new_n854), .A3(new_n1216), .ZN(new_n1217));
  OR4_X1    g1017(.A1(G387), .A2(new_n1215), .A3(G381), .A4(new_n1217), .ZN(G407));
  OAI211_X1 g1018(.A(G407), .B(G213), .C1(G343), .C2(new_n1215), .ZN(G409));
  INV_X1    g1019(.A(KEYINPUT61), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT60), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n705), .B1(new_n1221), .B2(new_n1191), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n1125), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1223), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1212), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n854), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1221), .A2(new_n1191), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n704), .A3(new_n1224), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(G384), .A3(new_n1212), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT125), .ZN(new_n1237));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(G343), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(G2897), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1235), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1240), .ZN(new_n1243));
  AOI211_X1 g1043(.A(KEYINPUT125), .B(new_n1243), .C1(new_n1228), .C2(new_n1234), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1237), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n704), .B(new_n1155), .C1(new_n1157), .C2(KEYINPUT120), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1131), .B(KEYINPUT57), .C1(new_n1133), .C2(new_n1152), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1188), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT123), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT123), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1159), .A2(new_n1250), .A3(G378), .A4(new_n1188), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1153), .A2(new_n1008), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1188), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1214), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1239), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1220), .B1(new_n1245), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1256), .B2(new_n1236), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1249), .A2(new_n1251), .B1(new_n1214), .B2(new_n1254), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(new_n1260), .A2(KEYINPUT62), .A3(new_n1239), .A4(new_n1235), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1257), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(new_n1216), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G387), .A2(new_n1077), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(G387), .A2(new_n1077), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(new_n1077), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1268), .A2(new_n1266), .A3(new_n1269), .A4(new_n1264), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1239), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1236), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1233), .B2(new_n1212), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n854), .B(new_n1211), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1241), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1243), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1235), .A2(new_n1241), .A3(new_n1240), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1237), .C1(new_n1239), .C2(new_n1260), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1279), .A2(new_n1220), .A3(new_n1274), .A4(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1276), .A4(new_n1236), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1256), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1236), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1262), .A2(new_n1274), .B1(new_n1287), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(G375), .A2(new_n1214), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1273), .A2(new_n1252), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1273), .B1(new_n1252), .B2(new_n1294), .ZN(new_n1296));
  OR3_X1    g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1235), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1235), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G402));
endmodule


