

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U561 ( .A(n732), .ZN(n706) );
  BUF_X1 U562 ( .A(n900), .Z(n527) );
  XNOR2_X1 U563 ( .A(n532), .B(n531), .ZN(n900) );
  NOR2_X1 U564 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U565 ( .A1(G8), .A2(n732), .ZN(n809) );
  NAND2_X1 U566 ( .A1(n686), .A2(n777), .ZN(n732) );
  NAND2_X1 U567 ( .A1(n900), .A2(G137), .ZN(n533) );
  NOR2_X1 U568 ( .A1(n809), .A2(n748), .ZN(n528) );
  XNOR2_X1 U569 ( .A(n695), .B(KEYINPUT93), .ZN(n696) );
  NOR2_X1 U570 ( .A1(G1966), .A2(n809), .ZN(n726) );
  NOR2_X1 U571 ( .A1(n743), .A2(n742), .ZN(n744) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n531) );
  AND2_X1 U573 ( .A1(n534), .A2(G2104), .ZN(n901) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n535) );
  NOR2_X1 U575 ( .A1(G651), .A2(n656), .ZN(n651) );
  XNOR2_X1 U576 ( .A(n536), .B(n535), .ZN(n537) );
  NOR2_X1 U577 ( .A1(n540), .A2(n539), .ZN(G160) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n905) );
  NAND2_X1 U579 ( .A1(G113), .A2(n905), .ZN(n530) );
  INV_X1 U580 ( .A(G2105), .ZN(n534) );
  NOR2_X1 U581 ( .A1(G2104), .A2(n534), .ZN(n906) );
  NAND2_X1 U582 ( .A1(G125), .A2(n906), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n540) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XNOR2_X1 U585 ( .A(n533), .B(KEYINPUT66), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G101), .A2(n901), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U588 ( .A1(G99), .A2(n901), .ZN(n547) );
  NAND2_X1 U589 ( .A1(G111), .A2(n905), .ZN(n542) );
  NAND2_X1 U590 ( .A1(G135), .A2(n527), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U592 ( .A1(n906), .A2(G123), .ZN(n543) );
  XOR2_X1 U593 ( .A(KEYINPUT18), .B(n543), .Z(n544) );
  NOR2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U595 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U596 ( .A(n548), .B(KEYINPUT76), .ZN(n1015) );
  XNOR2_X1 U597 ( .A(n1015), .B(G2096), .ZN(n549) );
  OR2_X1 U598 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G108), .ZN(G238) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n656) );
  NAND2_X1 U604 ( .A1(G52), .A2(n651), .ZN(n552) );
  INV_X1 U605 ( .A(G651), .ZN(n553) );
  NOR2_X1 U606 ( .A1(G543), .A2(n553), .ZN(n550) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(n550), .Z(n655) );
  NAND2_X1 U608 ( .A1(G64), .A2(n655), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n559) );
  NOR2_X1 U610 ( .A1(n656), .A2(n553), .ZN(n642) );
  NAND2_X1 U611 ( .A1(G77), .A2(n642), .ZN(n555) );
  NOR2_X1 U612 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U613 ( .A1(G90), .A2(n643), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n556), .Z(n557) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n557), .ZN(n558) );
  NOR2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G171) );
  INV_X1 U618 ( .A(G171), .ZN(G301) );
  NAND2_X1 U619 ( .A1(G138), .A2(n527), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G102), .A2(n901), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G114), .A2(n905), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G126), .A2(n906), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U625 ( .A1(n565), .A2(n564), .ZN(G164) );
  NAND2_X1 U626 ( .A1(G51), .A2(n651), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G63), .A2(n655), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U629 ( .A(KEYINPUT6), .B(n568), .ZN(n575) );
  NAND2_X1 U630 ( .A1(n643), .A2(G89), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G76), .A2(n642), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U634 ( .A(KEYINPUT5), .B(n572), .ZN(n573) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(n573), .ZN(n574) );
  NOR2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT7), .B(n576), .Z(G168) );
  NAND2_X1 U638 ( .A1(G94), .A2(G452), .ZN(n577) );
  XNOR2_X1 U639 ( .A(n577), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n841) );
  NAND2_X1 U643 ( .A1(n841), .A2(G567), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  XNOR2_X1 U645 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G81), .A2(n643), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT70), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G68), .A2(n642), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n655), .A2(G56), .ZN(n586) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n586), .Z(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n651), .A2(G43), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n935) );
  INV_X1 U657 ( .A(G860), .ZN(n617) );
  OR2_X1 U658 ( .A1(n935), .A2(n617), .ZN(G153) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U660 ( .A1(n651), .A2(G54), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G92), .A2(n643), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G66), .A2(n655), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n642), .A2(G79), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT72), .B(n593), .Z(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT15), .B(n598), .Z(n933) );
  INV_X1 U669 ( .A(G868), .ZN(n668) );
  NAND2_X1 U670 ( .A1(n933), .A2(n668), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G53), .A2(n651), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G65), .A2(n655), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G78), .A2(n642), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G91), .A2(n643), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n715) );
  INV_X1 U679 ( .A(n715), .ZN(G299) );
  XOR2_X1 U680 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT74), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n668), .A2(G286), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U685 ( .A(KEYINPUT75), .B(n610), .Z(G297) );
  NAND2_X1 U686 ( .A1(n617), .A2(G559), .ZN(n611) );
  INV_X1 U687 ( .A(n933), .ZN(n853) );
  NAND2_X1 U688 ( .A1(n611), .A2(n853), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n935), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G868), .A2(n853), .ZN(n613) );
  NOR2_X1 U692 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U694 ( .A1(G559), .A2(n853), .ZN(n616) );
  XOR2_X1 U695 ( .A(n935), .B(n616), .Z(n665) );
  NAND2_X1 U696 ( .A1(n617), .A2(n665), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G93), .A2(n643), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G67), .A2(n655), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G80), .A2(n642), .ZN(n620) );
  XNOR2_X1 U701 ( .A(KEYINPUT77), .B(n620), .ZN(n621) );
  NOR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n651), .A2(G55), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n667) );
  XNOR2_X1 U705 ( .A(n625), .B(n667), .ZN(G145) );
  NAND2_X1 U706 ( .A1(G73), .A2(n642), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT2), .B(n626), .Z(n629) );
  NAND2_X1 U708 ( .A1(n655), .A2(G61), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT78), .B(n627), .Z(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n643), .A2(G86), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n632), .B(KEYINPUT79), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G48), .A2(n651), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G47), .A2(n651), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G60), .A2(n655), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G72), .A2(n642), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G85), .A2(n643), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n641), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U724 ( .A1(G75), .A2(n642), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G88), .A2(n643), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G62), .A2(n655), .ZN(n646) );
  XNOR2_X1 U728 ( .A(n646), .B(KEYINPUT80), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n651), .A2(G50), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U731 ( .A1(n650), .A2(n649), .ZN(G166) );
  INV_X1 U732 ( .A(G166), .ZN(G303) );
  NAND2_X1 U733 ( .A1(G49), .A2(n651), .ZN(n653) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n656), .A2(G87), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(G288) );
  XOR2_X1 U739 ( .A(G305), .B(G290), .Z(n659) );
  XNOR2_X1 U740 ( .A(n667), .B(n659), .ZN(n660) );
  XOR2_X1 U741 ( .A(n660), .B(KEYINPUT19), .Z(n662) );
  XNOR2_X1 U742 ( .A(n715), .B(KEYINPUT81), .ZN(n661) );
  XNOR2_X1 U743 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n663), .B(G303), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n664), .B(G288), .ZN(n849) );
  XNOR2_X1 U746 ( .A(n665), .B(n849), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U748 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U759 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G96), .A2(n677), .ZN(n847) );
  NAND2_X1 U761 ( .A1(n847), .A2(G2106), .ZN(n683) );
  NAND2_X1 U762 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U763 ( .A1(G237), .A2(n678), .ZN(n679) );
  XOR2_X1 U764 ( .A(KEYINPUT82), .B(n679), .Z(n680) );
  NOR2_X1 U765 ( .A1(G238), .A2(n680), .ZN(n681) );
  XNOR2_X1 U766 ( .A(KEYINPUT83), .B(n681), .ZN(n848) );
  NAND2_X1 U767 ( .A1(n848), .A2(G567), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n922) );
  NOR2_X1 U769 ( .A1(n684), .A2(n922), .ZN(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT84), .ZN(n846) );
  NAND2_X1 U771 ( .A1(G36), .A2(n846), .ZN(G176) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n776) );
  INV_X1 U773 ( .A(n776), .ZN(n686) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NOR2_X1 U775 ( .A1(G2084), .A2(n732), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n728), .A2(n726), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n687), .A2(G8), .ZN(n688) );
  XNOR2_X1 U778 ( .A(n688), .B(KEYINPUT92), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n689), .B(KEYINPUT30), .ZN(n690) );
  NOR2_X1 U780 ( .A1(G168), .A2(n690), .ZN(n694) );
  NAND2_X1 U781 ( .A1(G1961), .A2(n732), .ZN(n692) );
  XOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .Z(n993) );
  NAND2_X1 U783 ( .A1(n706), .A2(n993), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n721) );
  AND2_X1 U785 ( .A1(G301), .A2(n721), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n697) );
  INV_X1 U787 ( .A(KEYINPUT31), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n697), .B(n696), .ZN(n725) );
  NAND2_X1 U789 ( .A1(n706), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U791 ( .A(G1956), .ZN(n965) );
  NOR2_X1 U792 ( .A1(n965), .A2(n706), .ZN(n699) );
  NOR2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n714) );
  NOR2_X1 U794 ( .A1(n715), .A2(n714), .ZN(n701) );
  XOR2_X1 U795 ( .A(n701), .B(KEYINPUT28), .Z(n719) );
  AND2_X1 U796 ( .A1(n706), .A2(G1996), .ZN(n702) );
  XOR2_X1 U797 ( .A(n702), .B(KEYINPUT26), .Z(n704) );
  NAND2_X1 U798 ( .A1(n732), .A2(G1341), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n935), .A2(n705), .ZN(n710) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n732), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G2067), .A2(n706), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n933), .A2(n711), .ZN(n709) );
  OR2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n933), .A2(n711), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U811 ( .A(n720), .B(KEYINPUT29), .ZN(n723) );
  NOR2_X1 U812 ( .A1(G301), .A2(n721), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n736) );
  NOR2_X1 U814 ( .A1(n726), .A2(n736), .ZN(n727) );
  XNOR2_X1 U815 ( .A(n727), .B(KEYINPUT94), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n728), .A2(G8), .ZN(n729) );
  NAND2_X1 U817 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U818 ( .A(KEYINPUT95), .B(n731), .ZN(n743) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n809), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U822 ( .A1(G303), .A2(n735), .ZN(n739) );
  INV_X1 U823 ( .A(n736), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G286), .A2(n737), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n740), .A2(G8), .ZN(n741) );
  XOR2_X1 U827 ( .A(KEYINPUT32), .B(n741), .Z(n742) );
  XNOR2_X1 U828 ( .A(n744), .B(KEYINPUT96), .ZN(n803) );
  INV_X1 U829 ( .A(n803), .ZN(n747) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n943), .A2(n745), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n940) );
  INV_X1 U835 ( .A(n940), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n528), .ZN(n751) );
  INV_X1 U837 ( .A(KEYINPUT64), .ZN(n750) );
  XNOR2_X1 U838 ( .A(n751), .B(n750), .ZN(n796) );
  INV_X1 U839 ( .A(KEYINPUT97), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n809), .A2(n753), .ZN(n794) );
  NAND2_X1 U841 ( .A1(n943), .A2(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n943), .A2(KEYINPUT97), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n809), .A2(n756), .ZN(n792) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n930) );
  NAND2_X1 U847 ( .A1(G105), .A2(n901), .ZN(n757) );
  XNOR2_X1 U848 ( .A(n757), .B(KEYINPUT38), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G117), .A2(n905), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G129), .A2(n906), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U852 ( .A(KEYINPUT88), .B(n760), .ZN(n763) );
  NAND2_X1 U853 ( .A1(G141), .A2(n527), .ZN(n761) );
  XNOR2_X1 U854 ( .A(KEYINPUT89), .B(n761), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n920) );
  NAND2_X1 U857 ( .A1(G1996), .A2(n920), .ZN(n766) );
  XOR2_X1 U858 ( .A(KEYINPUT90), .B(n766), .Z(n774) );
  NAND2_X1 U859 ( .A1(G131), .A2(n527), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G95), .A2(n901), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G107), .A2(n905), .ZN(n770) );
  NAND2_X1 U863 ( .A1(G119), .A2(n906), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n897) );
  AND2_X1 U866 ( .A1(n897), .A2(G1991), .ZN(n773) );
  NOR2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n814) );
  XNOR2_X1 U868 ( .A(KEYINPUT85), .B(G1986), .ZN(n775) );
  XNOR2_X1 U869 ( .A(n775), .B(G290), .ZN(n950) );
  NAND2_X1 U870 ( .A1(n814), .A2(n950), .ZN(n778) );
  NOR2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n820) );
  NAND2_X1 U872 ( .A1(n778), .A2(n820), .ZN(n811) );
  AND2_X1 U873 ( .A1(n930), .A2(n811), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n779) );
  XNOR2_X1 U875 ( .A(n779), .B(KEYINPUT86), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G140), .A2(n527), .ZN(n781) );
  NAND2_X1 U877 ( .A1(G104), .A2(n901), .ZN(n780) );
  NAND2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G116), .A2(n905), .ZN(n784) );
  NAND2_X1 U881 ( .A1(G128), .A2(n906), .ZN(n783) );
  NAND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U883 ( .A(n785), .B(KEYINPUT35), .Z(n786) );
  NOR2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U885 ( .A(n789), .B(n788), .ZN(n915) );
  XOR2_X1 U886 ( .A(KEYINPUT37), .B(G2067), .Z(n819) );
  AND2_X1 U887 ( .A1(n915), .A2(n819), .ZN(n1025) );
  NAND2_X1 U888 ( .A1(n1025), .A2(n820), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n790), .A2(n800), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n797) );
  INV_X1 U891 ( .A(n797), .ZN(n793) );
  NOR2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n797), .A2(KEYINPUT33), .ZN(n798) );
  AND2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n830) );
  INV_X1 U896 ( .A(n800), .ZN(n828) );
  NAND2_X1 U897 ( .A1(G166), .A2(G8), .ZN(n801) );
  NOR2_X1 U898 ( .A1(G2090), .A2(n801), .ZN(n802) );
  OR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n805) );
  AND2_X1 U900 ( .A1(n809), .A2(n811), .ZN(n804) );
  AND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n826) );
  NOR2_X1 U902 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XNOR2_X1 U903 ( .A(n806), .B(KEYINPUT24), .ZN(n807) );
  XNOR2_X1 U904 ( .A(KEYINPUT91), .B(n807), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n824) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n920), .ZN(n1020) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n897), .ZN(n1013) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n812) );
  XNOR2_X1 U910 ( .A(KEYINPUT98), .B(n812), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n1013), .A2(n813), .ZN(n815) );
  INV_X1 U912 ( .A(n814), .ZN(n1017) );
  NOR2_X1 U913 ( .A1(n815), .A2(n1017), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n1020), .A2(n816), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT39), .B(n817), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n818), .A2(n820), .ZN(n822) );
  NOR2_X1 U917 ( .A1(n819), .A2(n915), .ZN(n1034) );
  NAND2_X1 U918 ( .A1(n1034), .A2(n820), .ZN(n821) );
  AND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  OR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U924 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U925 ( .A(G1348), .B(G2454), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n832), .B(G2430), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(G1341), .ZN(n839) );
  XOR2_X1 U928 ( .A(G2443), .B(G2427), .Z(n835) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U931 ( .A(G2451), .B(G2435), .Z(n836) );
  XNOR2_X1 U932 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n840), .A2(G14), .ZN(n925) );
  XNOR2_X1 U935 ( .A(KEYINPUT99), .B(n925), .ZN(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n841), .ZN(G217) );
  INV_X1 U937 ( .A(G661), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G2), .A2(G15), .ZN(n842) );
  NOR2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT100), .B(n844), .Z(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U944 ( .A(G120), .ZN(G236) );
  INV_X1 U945 ( .A(G96), .ZN(G221) );
  INV_X1 U946 ( .A(G69), .ZN(G235) );
  NOR2_X1 U947 ( .A1(n848), .A2(n847), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  XOR2_X1 U949 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n851) );
  XNOR2_X1 U950 ( .A(G171), .B(n849), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U952 ( .A(G286), .B(n852), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n935), .B(n853), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  NOR2_X1 U955 ( .A1(G37), .A2(n856), .ZN(G397) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2090), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT42), .ZN(n867) );
  XOR2_X1 U958 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT103), .B(G2096), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(G2100), .B(G2072), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(G2678), .B(KEYINPUT43), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(G227) );
  XOR2_X1 U968 ( .A(G1986), .B(G1971), .Z(n869) );
  XNOR2_X1 U969 ( .A(G1961), .B(G1956), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(n870), .B(G2474), .Z(n872) );
  XNOR2_X1 U972 ( .A(G1996), .B(G1991), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U974 ( .A(KEYINPUT41), .B(G1976), .Z(n874) );
  XNOR2_X1 U975 ( .A(G1966), .B(G1981), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U978 ( .A1(G124), .A2(n906), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n877), .B(KEYINPUT44), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(KEYINPUT104), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G112), .A2(n905), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G136), .A2(n527), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G100), .A2(n901), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(G162) );
  XOR2_X1 U987 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT108), .B(KEYINPUT48), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G139), .A2(n527), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G103), .A2(n901), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n905), .A2(G115), .ZN(n889) );
  XNOR2_X1 U994 ( .A(KEYINPUT107), .B(n889), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n906), .A2(G127), .ZN(n890) );
  XOR2_X1 U996 ( .A(KEYINPUT106), .B(n890), .Z(n891) );
  NOR2_X1 U997 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U998 ( .A(n893), .B(KEYINPUT47), .ZN(n894) );
  NOR2_X1 U999 ( .A1(n895), .A2(n894), .ZN(n1027) );
  XOR2_X1 U1000 ( .A(n896), .B(n1027), .Z(n899) );
  XOR2_X1 U1001 ( .A(G160), .B(n897), .Z(n898) );
  XNOR2_X1 U1002 ( .A(n899), .B(n898), .ZN(n914) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n527), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(G106), .A2(n901), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1006 ( .A(n904), .B(KEYINPUT45), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(G118), .A2(n905), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(G130), .A2(n906), .ZN(n907) );
  NAND2_X1 U1009 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(KEYINPUT105), .B(n909), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n912), .B(G162), .ZN(n913) );
  XOR2_X1 U1013 ( .A(n914), .B(n913), .Z(n917) );
  XOR2_X1 U1014 ( .A(n915), .B(G164), .Z(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1016 ( .A(n1015), .B(n918), .Z(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n921), .ZN(G395) );
  INV_X1 U1019 ( .A(n922), .ZN(G319) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n924), .ZN(n929) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n925), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT112), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(G395), .A2(n927), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1028 ( .A(G16), .B(KEYINPUT56), .ZN(n955) );
  XNOR2_X1 U1029 ( .A(G1966), .B(G168), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT57), .B(n932), .ZN(n953) );
  XNOR2_X1 U1032 ( .A(G1348), .B(KEYINPUT118), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(n933), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(G1341), .B(n935), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(G301), .B(G1961), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G299), .B(G1956), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n948) );
  XOR2_X1 U1042 ( .A(G1971), .B(G303), .Z(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n946), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT120), .B(n951), .Z(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n986) );
  INV_X1 U1049 ( .A(G16), .ZN(n984) );
  XNOR2_X1 U1050 ( .A(G1986), .B(KEYINPUT126), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(G24), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT124), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n960), .B(KEYINPUT125), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1058 ( .A(KEYINPUT58), .B(n963), .Z(n981) );
  XOR2_X1 U1059 ( .A(G1961), .B(G5), .Z(n976) );
  XOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .Z(n964) );
  XNOR2_X1 U1061 ( .A(G4), .B(n964), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(G20), .B(n965), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(n966), .B(KEYINPUT121), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G6), .B(G1981), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1068 ( .A(KEYINPUT122), .B(n971), .Z(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n974), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G21), .B(G1966), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT123), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT61), .B(n982), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n1009) );
  XNOR2_X1 U1079 ( .A(KEYINPUT116), .B(G2084), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(KEYINPUT54), .B(G34), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n987), .B(KEYINPUT115), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n989), .B(n988), .ZN(n1004) );
  XNOR2_X1 U1083 ( .A(G2090), .B(G35), .ZN(n1002) );
  XOR2_X1 U1084 ( .A(G25), .B(G1991), .Z(n990) );
  NAND2_X1 U1085 ( .A1(n990), .A2(G28), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1996), .B(G32), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(G33), .B(G2072), .ZN(n991) );
  NOR2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(G2067), .B(G26), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(G27), .B(n993), .ZN(n994) );
  NOR2_X1 U1091 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(KEYINPUT53), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1097 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n1005) );
  XNOR2_X1 U1098 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(G29), .A2(n1007), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(G11), .A2(n1010), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(KEYINPUT127), .ZN(n1040) );
  XOR2_X1 U1103 ( .A(G2084), .B(G160), .Z(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(G2090), .B(G162), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(n1018), .B(KEYINPUT113), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1110 ( .A(KEYINPUT51), .B(n1021), .Z(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT114), .B(n1026), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(G2072), .B(n1027), .Z(n1029) );
  XOR2_X1 U1115 ( .A(G164), .B(G2078), .Z(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1117 ( .A(KEYINPUT50), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(KEYINPUT52), .B(n1035), .ZN(n1037) );
  INV_X1 U1121 ( .A(KEYINPUT55), .ZN(n1036) );
  NAND2_X1 U1122 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(G29), .ZN(n1039) );
  NAND2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

