//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT78), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  AOI21_X1  g004(.A(G107), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT80), .B1(new_n192), .B2(G104), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n187), .A3(G107), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n191), .B2(new_n196), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n187), .A2(KEYINPUT3), .A3(G107), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n191), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n188), .A2(new_n190), .A3(G107), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n197), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G113), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G116), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n207), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n220), .B2(new_n208), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT2), .B(G113), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n218), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n206), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n216), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n222), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n224), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT67), .A4(new_n222), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n189), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n187), .A2(KEYINPUT78), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n192), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n198), .B1(new_n234), .B2(KEYINPUT3), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n203), .B1(new_n235), .B2(new_n202), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT4), .B1(new_n201), .B2(new_n204), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n230), .B(new_n231), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n202), .B(new_n199), .C1(new_n191), .C2(new_n200), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n225), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n225), .B(new_n246), .C1(new_n238), .C2(new_n244), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n251), .A3(new_n247), .ZN(new_n252));
  INV_X1    g066(.A(G224), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G953), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n258), .A3(G146), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G143), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n256), .A2(new_n258), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(new_n261), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n264), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT64), .B(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(G146), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT1), .B1(new_n255), .B2(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n262), .A2(new_n279), .A3(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(G128), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n262), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n275), .B2(G146), .ZN(new_n283));
  INV_X1    g097(.A(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT1), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n276), .A2(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n271), .A2(new_n272), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n254), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n290), .ZN(new_n292));
  INV_X1    g106(.A(new_n254), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n288), .A4(new_n273), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n250), .A2(new_n252), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n221), .A2(new_n205), .A3(new_n224), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n246), .B(KEYINPUT8), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n218), .A2(KEYINPUT5), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n212), .A2(new_n299), .B1(new_n223), .B2(new_n218), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n298), .C1(new_n205), .C2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n249), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT7), .B(new_n293), .C1(new_n289), .C2(new_n290), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n292), .A2(new_n288), .A3(new_n273), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT88), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n310), .B(KEYINPUT87), .Z(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n296), .A2(new_n307), .A3(new_n310), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n311), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n296), .B2(new_n307), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(new_n309), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G214), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT69), .B(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n284), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n209), .A2(G128), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n326), .B1(KEYINPUT73), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT73), .B(KEYINPUT23), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n332), .B(new_n327), .C1(new_n333), .C2(new_n326), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n330), .B1(new_n334), .B2(G110), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n287), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n339), .A2(KEYINPUT76), .A3(G146), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT76), .B1(new_n339), .B2(G146), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT75), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT16), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n336), .A4(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n348), .A2(new_n351), .A3(G146), .A4(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n261), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n353), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n328), .A2(new_n329), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n328), .B2(new_n329), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n358), .A2(new_n359), .B1(new_n334), .B2(G110), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n343), .A2(new_n353), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n325), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n360), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n335), .A2(new_n342), .A3(new_n353), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n362), .A3(new_n365), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(new_n369), .B2(new_n325), .ZN(new_n370));
  INV_X1    g184(.A(G902), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT25), .A3(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n364), .A2(new_n362), .A3(new_n365), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n325), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n325), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(G234), .B2(new_n371), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(G902), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n370), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G237), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n322), .A2(G210), .A3(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT26), .B(G101), .Z(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n281), .A2(new_n276), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n283), .A2(new_n285), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT11), .ZN(new_n396));
  INV_X1    g210(.A(G134), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(G137), .ZN(new_n398));
  INV_X1    g212(.A(G137), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT11), .A3(G134), .ZN(new_n400));
  INV_X1    g214(.A(G131), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(G137), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n397), .A2(G137), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n399), .A2(G134), .ZN(new_n405));
  OAI21_X1  g219(.A(G131), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n394), .A2(new_n395), .B1(KEYINPUT68), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n276), .A2(new_n268), .B1(new_n283), .B2(new_n260), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G131), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n408), .A2(new_n410), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT28), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n230), .A2(new_n231), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n407), .A2(KEYINPUT68), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n284), .B1(new_n277), .B2(KEYINPUT65), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n257), .A2(G143), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n261), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n280), .A2(new_n420), .B1(new_n423), .B2(new_n274), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n259), .A2(new_n262), .A3(new_n285), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n419), .B(new_n410), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n411), .A2(new_n414), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT28), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n417), .ZN(new_n431));
  INV_X1    g245(.A(new_n414), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n270), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n407), .B1(new_n394), .B2(new_n395), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n393), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n428), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n427), .B(new_n439), .C1(new_n286), .C2(new_n407), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n415), .B2(new_n439), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n438), .B1(new_n441), .B2(new_n431), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT31), .B1(new_n442), .B2(new_n393), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT30), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n426), .B2(new_n427), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n431), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(KEYINPUT31), .A3(new_n428), .A4(new_n393), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n437), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n450));
  NOR2_X1   g264(.A1(G472), .A2(G902), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n446), .A2(new_n428), .A3(new_n393), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT31), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n436), .B1(new_n455), .B2(new_n447), .ZN(new_n456));
  INV_X1    g270(.A(new_n451), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT32), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n430), .A2(new_n435), .A3(new_n393), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT71), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n446), .A2(new_n428), .ZN(new_n462));
  INV_X1    g276(.A(new_n393), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n430), .A2(new_n465), .A3(new_n435), .A4(new_n393), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n426), .A2(new_n427), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n431), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n429), .B2(new_n418), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n393), .A2(KEYINPUT29), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G472), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n387), .B1(new_n459), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G116), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n213), .A2(G122), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n192), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT14), .B1(new_n477), .B2(G116), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n213), .A3(G122), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT95), .A4(new_n478), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n482), .B1(new_n493), .B2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n256), .A2(new_n258), .A3(G128), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT92), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n256), .A2(new_n258), .A3(new_n497), .A4(G128), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n255), .A2(G128), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT93), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n503), .B(new_n500), .C1(new_n496), .C2(new_n498), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n502), .A2(new_n504), .A3(new_n397), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n497), .B1(new_n275), .B2(G128), .ZN(new_n506));
  AND4_X1   g320(.A1(new_n497), .A2(new_n256), .A3(new_n258), .A4(G128), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n503), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n499), .A2(KEYINPUT93), .A3(new_n501), .ZN(new_n510));
  AOI21_X1  g324(.A(G134), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n494), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n499), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n501), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n499), .A2(new_n513), .ZN(new_n516));
  OAI21_X1  g330(.A(G134), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n397), .B1(new_n502), .B2(new_n504), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n480), .B(new_n192), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT9), .B(G234), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n521), .A2(new_n382), .A3(G953), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n512), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n512), .B2(new_n520), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n371), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT96), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT96), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(new_n371), .C1(new_n523), .C2(new_n524), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n528), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n371), .B(new_n532), .C1(new_n523), .C2(new_n524), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(KEYINPUT97), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(KEYINPUT97), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G953), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT69), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n538), .A2(new_n540), .A3(G214), .A4(new_n388), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n275), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n322), .A2(G143), .A3(G214), .A4(new_n388), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G131), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n401), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(KEYINPUT17), .A3(G131), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n550), .A2(new_n355), .A3(new_n353), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n545), .A2(new_n552), .A3(new_n546), .A4(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n339), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n342), .B1(new_n261), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT18), .A2(G131), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n542), .A2(new_n543), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n544), .A2(KEYINPUT18), .A3(G131), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(G113), .B(G122), .Z(new_n561));
  XOR2_X1   g375(.A(KEYINPUT89), .B(G104), .Z(new_n562));
  XOR2_X1   g376(.A(new_n561), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT90), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n554), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n545), .A2(new_n547), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT19), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n339), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n261), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n353), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n560), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n563), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(G475), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT20), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(new_n565), .ZN(new_n579));
  INV_X1    g393(.A(new_n563), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n554), .B2(new_n560), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n371), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n576), .A2(new_n578), .B1(new_n582), .B2(G475), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n537), .A2(G952), .ZN(new_n585));
  INV_X1    g399(.A(G234), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n388), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n371), .B(new_n322), .C1(G234), .C2(G237), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT21), .B(G898), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n536), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G221), .B1(new_n521), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n371), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT78), .B(G104), .ZN(new_n597));
  AOI21_X1  g411(.A(G101), .B1(new_n597), .B2(G107), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n598), .B(new_n199), .C1(new_n200), .C2(new_n191), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT1), .B1(new_n275), .B2(G146), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(G128), .B1(new_n262), .B2(new_n259), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n599), .B(new_n197), .C1(new_n601), .C2(new_n425), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n205), .A2(new_n286), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n414), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT84), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n604), .A2(new_n611), .A3(new_n607), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n611), .B1(new_n604), .B2(new_n607), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n612), .B(new_n606), .C1(new_n602), .C2(new_n603), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT84), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n394), .B2(new_n395), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n602), .A2(new_n620), .B1(new_n206), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n239), .A2(G101), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n599), .A3(KEYINPUT4), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n624), .B(new_n411), .C1(new_n242), .C2(new_n243), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n432), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n322), .A2(G227), .ZN(new_n627));
  XOR2_X1   g441(.A(G110), .B(G140), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n616), .A2(new_n619), .A3(new_n626), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n626), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n432), .B1(new_n622), .B2(new_n625), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n596), .B1(new_n635), .B2(new_n595), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n626), .B1(new_n618), .B2(new_n617), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT82), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n626), .B(KEYINPUT82), .C1(new_n618), .C2(new_n617), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n629), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT83), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n632), .B2(new_n629), .ZN(new_n643));
  INV_X1    g457(.A(new_n633), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n626), .A2(KEYINPUT83), .A3(new_n630), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n646), .A3(G469), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n594), .B1(new_n636), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n321), .A2(new_n476), .A3(new_n592), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT98), .B(G101), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT99), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(G3));
  AND3_X1   g466(.A1(new_n296), .A2(new_n307), .A3(new_n310), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n310), .B1(new_n296), .B2(new_n307), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n319), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT100), .ZN(new_n656));
  INV_X1    g470(.A(new_n591), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n319), .C1(new_n653), .C2(new_n654), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n631), .A2(new_n634), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n595), .A3(new_n371), .ZN(new_n663));
  INV_X1    g477(.A(new_n596), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n647), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n593), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n456), .B2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n449), .A2(new_n451), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n666), .A2(new_n387), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n512), .A2(new_n520), .A3(new_n522), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n512), .A2(new_n520), .ZN(new_n674));
  INV_X1    g488(.A(new_n522), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n512), .A2(new_n520), .A3(KEYINPUT102), .A4(new_n522), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n676), .A3(KEYINPUT33), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT101), .B(KEYINPUT33), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n523), .B2(new_n524), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n527), .A2(G902), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n678), .A2(KEYINPUT103), .A3(new_n680), .A4(new_n681), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n584), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n661), .A2(new_n670), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n187), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  NAND2_X1  g507(.A1(new_n582), .A2(G475), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n695), .B(new_n577), .C1(new_n573), .C2(new_n574), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n577), .B1(new_n573), .B2(new_n574), .ZN(new_n697));
  INV_X1    g511(.A(new_n574), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT20), .B(new_n698), .C1(new_n565), .C2(new_n572), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n696), .B1(new_n700), .B2(new_n695), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n536), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n661), .A2(new_n670), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT35), .B(G107), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G9));
  INV_X1    g519(.A(new_n383), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n372), .B2(new_n380), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n376), .A2(KEYINPUT36), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n366), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n385), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n666), .A2(new_n669), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n321), .A3(new_n592), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT37), .B(G110), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G12));
  INV_X1    g530(.A(new_n310), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n308), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n313), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n658), .B1(new_n719), .B2(new_n319), .ZN(new_n720));
  INV_X1    g534(.A(new_n659), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n589), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n587), .B1(new_n723), .B2(G900), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n536), .A2(new_n694), .A3(new_n701), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n712), .B1(new_n459), .B2(new_n475), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n648), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G128), .ZN(G30));
  OAI21_X1  g542(.A(KEYINPUT38), .B1(new_n314), .B2(new_n317), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n316), .A2(new_n309), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT38), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n313), .A4(new_n312), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n442), .A2(new_n463), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n463), .A2(new_n428), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n371), .B1(new_n735), .B2(new_n470), .ZN(new_n736));
  OAI21_X1  g550(.A(G472), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n456), .A2(KEYINPUT32), .A3(new_n457), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT97), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n533), .B(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n583), .B1(new_n742), .B2(new_n531), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n384), .A2(new_n710), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n320), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n733), .A2(new_n740), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT40), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n724), .B(KEYINPUT39), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT106), .B1(new_n648), .B2(new_n748), .ZN(new_n749));
  AND4_X1   g563(.A1(KEYINPUT106), .A2(new_n665), .A3(new_n593), .A4(new_n748), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  INV_X1    g566(.A(new_n748), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n666), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n648), .A2(KEYINPUT106), .A3(new_n748), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(KEYINPUT40), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n746), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n275), .ZN(G45));
  AND3_X1   g572(.A1(new_n687), .A2(new_n584), .A3(new_n724), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n722), .A2(new_n759), .A3(new_n648), .A4(new_n726), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT107), .B(G146), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G48));
  NAND2_X1  g576(.A1(new_n459), .A2(new_n475), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n707), .B1(new_n370), .B2(new_n385), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n635), .A2(new_n595), .ZN(new_n765));
  AOI211_X1 g579(.A(G469), .B(G902), .C1(new_n631), .C2(new_n634), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n765), .A2(new_n766), .A3(new_n594), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n660), .A3(new_n688), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT41), .B(G113), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G15));
  NAND4_X1  g585(.A1(new_n702), .A2(new_n657), .A3(new_n659), .A4(new_n656), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT108), .B1(new_n772), .B2(new_n768), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n774), .A2(new_n661), .A3(new_n775), .A4(new_n702), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G116), .ZN(G18));
  NAND2_X1  g592(.A1(new_n726), .A2(new_n592), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n767), .A2(new_n656), .A3(new_n659), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n209), .ZN(G21));
  NAND2_X1  g596(.A1(new_n455), .A2(new_n447), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n471), .A2(new_n393), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n457), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n449), .A2(new_n371), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(G472), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n767), .A2(new_n764), .A3(new_n657), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n656), .A2(new_n743), .A3(new_n659), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n477), .ZN(G24));
  AND2_X1   g605(.A1(new_n744), .A2(new_n787), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n722), .A2(new_n759), .A3(new_n767), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G125), .ZN(G27));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n314), .A2(new_n317), .A3(new_n320), .A4(new_n594), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n647), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n641), .A2(new_n646), .A3(KEYINPUT109), .A4(G469), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n636), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n476), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n759), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n795), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n459), .A2(new_n804), .B1(G472), .B2(new_n474), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n452), .A2(new_n458), .A3(KEYINPUT110), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n387), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n653), .B1(new_n309), .B2(new_n316), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n319), .A3(new_n730), .A4(new_n593), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n798), .A2(new_n636), .A3(new_n799), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(KEYINPUT42), .A3(new_n759), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n803), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  NAND4_X1  g628(.A1(new_n476), .A2(new_n725), .A3(new_n796), .A4(new_n800), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G134), .ZN(G36));
  NOR2_X1   g630(.A1(new_n753), .A2(new_n594), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n641), .A2(new_n646), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n641), .A2(new_n646), .A3(KEYINPUT45), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(G469), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n664), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT46), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n766), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n664), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n818), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n457), .B1(new_n783), .B2(new_n437), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n786), .B2(G472), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT111), .B1(new_n830), .B2(new_n712), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n744), .A2(new_n669), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n687), .A2(new_n583), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT43), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT43), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n687), .A2(new_n837), .A3(new_n583), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(KEYINPUT44), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n314), .A2(new_n320), .A3(new_n317), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n828), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT44), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n838), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n830), .A2(new_n712), .A3(KEYINPUT111), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n832), .B1(new_n744), .B2(new_n669), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n842), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT112), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n834), .A2(new_n836), .A3(new_n838), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n842), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n841), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(new_n399), .ZN(G39));
  NAND2_X1  g667(.A1(new_n824), .A2(new_n825), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n663), .A3(new_n827), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n593), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT47), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT47), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n858), .A3(new_n593), .ZN(new_n859));
  INV_X1    g673(.A(new_n840), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n802), .A2(new_n860), .A3(new_n763), .A4(new_n764), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(G140), .ZN(G42));
  NAND3_X1  g677(.A1(new_n764), .A2(new_n588), .A3(new_n787), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n843), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n767), .A2(new_n320), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n767), .A2(KEYINPUT115), .A3(new_n320), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n733), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n870), .A3(KEYINPUT50), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n765), .A2(new_n766), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n796), .A2(new_n588), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n843), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n792), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n857), .A2(new_n859), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n594), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n840), .A3(new_n865), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n764), .A2(new_n459), .A3(new_n737), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n877), .A2(KEYINPUT116), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT116), .B1(new_n877), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n687), .A2(new_n584), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n880), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT51), .A4(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n878), .A2(new_n807), .ZN(new_n894));
  NAND2_X1  g708(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n895));
  OR2_X1    g709(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n585), .C1(new_n894), .C2(new_n895), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n886), .A2(new_n689), .A3(new_n887), .ZN(new_n899));
  INV_X1    g713(.A(new_n780), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n865), .A2(KEYINPUT117), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT117), .B1(new_n865), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n893), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n769), .A2(new_n781), .A3(new_n790), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n813), .A3(new_n777), .ZN(new_n907));
  INV_X1    g721(.A(new_n536), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n688), .B1(new_n908), .B2(new_n584), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n319), .B(new_n657), .C1(new_n314), .C2(new_n317), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n670), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n714), .A3(new_n649), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n759), .A2(new_n792), .A3(new_n796), .A4(new_n800), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n694), .A2(new_n724), .ZN(new_n915));
  AND4_X1   g729(.A1(new_n531), .A2(new_n701), .A3(new_n742), .A4(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n726), .A2(new_n916), .A3(new_n648), .A4(new_n840), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n815), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n907), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n724), .A2(new_n593), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n707), .A2(new_n711), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n740), .A2(new_n800), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n656), .A2(new_n743), .A3(new_n659), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n760), .A2(new_n793), .A3(new_n925), .A4(new_n727), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT52), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n720), .A2(new_n666), .A3(new_n721), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n928), .B(new_n726), .C1(new_n725), .C2(new_n759), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT52), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n929), .A2(new_n930), .A3(new_n793), .A4(new_n925), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n920), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n913), .A2(new_n918), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(new_n777), .A3(new_n813), .A4(new_n906), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n927), .A2(new_n931), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT53), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT54), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT114), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n907), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n913), .A2(new_n918), .A3(new_n937), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n906), .A2(new_n813), .A3(new_n777), .A4(KEYINPUT114), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n941), .A2(new_n932), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n905), .A2(new_n948), .B1(G952), .B2(G953), .ZN(new_n949));
  INV_X1    g763(.A(new_n835), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n387), .A2(new_n320), .A3(new_n594), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT49), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n876), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT113), .Z(new_n954));
  INV_X1    g768(.A(new_n733), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n740), .B1(new_n952), .B2(new_n876), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n957), .ZN(G75));
  NOR2_X1   g772(.A1(new_n322), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n371), .B1(new_n944), .B2(new_n946), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(new_n311), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n250), .A2(new_n252), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT119), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n295), .B(KEYINPUT55), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT56), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n960), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n961), .A2(G210), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n970), .B2(new_n967), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(G51));
  XNOR2_X1  g786(.A(new_n596), .B(KEYINPUT57), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n662), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n961), .A2(G469), .A3(new_n822), .A4(new_n821), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n959), .B1(new_n977), .B2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n961), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n573), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n959), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT120), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n961), .A2(new_n984), .A3(new_n573), .A4(new_n980), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n961), .A2(new_n573), .A3(new_n980), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT120), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(G60));
  AND2_X1   g802(.A1(new_n678), .A2(new_n680), .ZN(new_n989));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT59), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n989), .B(new_n991), .C1(new_n974), .C2(new_n975), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n960), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n989), .B1(new_n948), .B2(new_n991), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(G63));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  NAND2_X1  g810(.A1(G217), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT60), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n944), .B2(new_n946), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n709), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n960), .B1(new_n999), .B2(new_n370), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n370), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n944), .A2(new_n946), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n998), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1006), .A2(KEYINPUT61), .A3(new_n960), .A4(new_n1000), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(G66));
  INV_X1    g822(.A(new_n590), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n537), .B1(new_n1009), .B2(G224), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n906), .A2(new_n777), .ZN(new_n1011));
  INV_X1    g825(.A(new_n913), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n1013), .B2(new_n322), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n964), .B1(G898), .B2(new_n322), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT121), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1014), .B(new_n1016), .ZN(G69));
  INV_X1    g831(.A(new_n322), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n441), .B(KEYINPUT122), .Z(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(new_n568), .ZN(new_n1020));
  OAI211_X1 g834(.A(G900), .B(new_n1018), .C1(new_n1020), .C2(G227), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(G227), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT124), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n754), .A2(new_n755), .ZN(new_n1024));
  INV_X1    g838(.A(new_n909), .ZN(new_n1025));
  INV_X1    g839(.A(new_n476), .ZN(new_n1026));
  NOR4_X1   g840(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n860), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1023), .B1(new_n852), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1027), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n849), .A2(new_n850), .A3(new_n842), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n850), .B1(new_n849), .B2(new_n842), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g846(.A(KEYINPUT124), .B(new_n1029), .C1(new_n1032), .C2(new_n841), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n760), .A2(new_n793), .A3(new_n727), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT62), .B1(new_n757), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n862), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n751), .A2(new_n756), .ZN(new_n1038));
  INV_X1    g852(.A(new_n746), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n760), .A2(new_n793), .A3(new_n727), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT62), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT123), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT123), .A4(new_n1042), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1037), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n1034), .A2(new_n1047), .ZN(new_n1048));
  OR2_X1    g862(.A1(new_n1048), .A2(new_n1020), .ZN(new_n1049));
  AND3_X1   g863(.A1(new_n929), .A2(new_n793), .A3(new_n815), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n828), .A2(new_n924), .A3(new_n807), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n862), .A2(new_n1050), .A3(new_n813), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1052), .A2(new_n852), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1018), .B1(new_n1053), .B2(new_n1020), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1022), .B1(new_n1049), .B2(new_n1054), .ZN(G72));
  XNOR2_X1  g869(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1056));
  NAND2_X1  g870(.A1(G472), .A2(G902), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g873(.A(new_n453), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n442), .A2(new_n393), .ZN(new_n1061));
  XNOR2_X1  g875(.A(new_n1061), .B(KEYINPUT127), .ZN(new_n1062));
  OAI221_X1 g876(.A(new_n1059), .B1(new_n1060), .B2(new_n1062), .C1(new_n933), .C2(new_n938), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n735), .B1(new_n431), .B2(new_n441), .ZN(new_n1064));
  NOR3_X1   g878(.A1(new_n1013), .A2(new_n1052), .A3(new_n852), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1064), .B1(new_n1065), .B2(new_n1058), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1063), .A2(new_n960), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g881(.A(new_n1013), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1034), .A2(new_n1047), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1069), .A2(KEYINPUT126), .A3(new_n1059), .ZN(new_n1070));
  AND2_X1   g884(.A1(new_n1070), .A2(new_n734), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1069), .A2(new_n1059), .ZN(new_n1072));
  INV_X1    g886(.A(KEYINPUT126), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1067), .B1(new_n1071), .B2(new_n1074), .ZN(G57));
endmodule


