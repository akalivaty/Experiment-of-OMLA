//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G250), .B1(G257), .B2(G264), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n201), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n216), .A2(G50), .A3(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n214), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT65), .Z(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  INV_X1    g0027(.A(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G116), .ZN(new_n229));
  INV_X1    g0029(.A(G270), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n202), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n232));
  INV_X1    g0032(.A(G77), .ZN(new_n233));
  INV_X1    g0033(.A(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G264), .ZN(new_n235));
  OAI221_X1 g0035(.A(new_n232), .B1(new_n233), .B2(new_n234), .C1(new_n206), .C2(new_n235), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n209), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n226), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT2), .B(G226), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n256), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n220), .B1(new_n209), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n202), .B1(new_n256), .B2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n202), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n264), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT8), .B(G58), .Z(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT69), .B1(new_n263), .B2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(new_n221), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n271), .A2(new_n275), .B1(G150), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT70), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n277), .A2(new_n278), .B1(G20), .B2(new_n203), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n269), .B1(new_n281), .B2(KEYINPUT71), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n281), .A2(KEYINPUT71), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n256), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  INV_X1    g0091(.A(new_n220), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n220), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n302), .B2(new_n228), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT3), .B(G33), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(G222), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(G1698), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT68), .B(G223), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(new_n233), .B2(new_n304), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n303), .B1(new_n297), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G169), .B2(new_n310), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n285), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(G190), .B2(new_n310), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n283), .A2(KEYINPUT9), .A3(new_n284), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  INV_X1    g0119(.A(new_n284), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n282), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n317), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT10), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(new_n317), .C1(new_n318), .C2(new_n321), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n314), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n261), .A2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT74), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n265), .B(G77), .C1(G1), .C2(new_n221), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n271), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT15), .B(G87), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n275), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n328), .B(new_n329), .C1(new_n270), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n297), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n304), .A2(G232), .A3(new_n305), .ZN(new_n337));
  XOR2_X1   g0137(.A(new_n337), .B(KEYINPUT73), .Z(new_n338));
  INV_X1    g0138(.A(G238), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n307), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(G107), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n336), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n295), .B1(new_n302), .B2(new_n234), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n335), .B1(new_n348), .B2(G190), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n315), .B2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n311), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n346), .B2(new_n347), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n335), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G274), .B1(new_n296), .B2(new_n220), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n288), .B2(new_n289), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G238), .B2(new_n301), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  INV_X1    g0160(.A(G232), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G1698), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G226), .B2(G1698), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(new_n344), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n297), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n358), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G200), .B2(new_n368), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT77), .ZN(new_n372));
  INV_X1    g0172(.A(G68), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n262), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n265), .B(G68), .C1(G1), .C2(new_n221), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n275), .A2(G77), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n221), .A2(G68), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n233), .B1(new_n272), .B2(new_n274), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT75), .B1(new_n383), .B2(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n276), .A2(G50), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n264), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT76), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(KEYINPUT76), .A3(new_n264), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n377), .B1(new_n391), .B2(KEYINPUT11), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT11), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n372), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n386), .A2(KEYINPUT76), .A3(new_n264), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT76), .B1(new_n386), .B2(new_n264), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT11), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n375), .A2(new_n376), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n394), .A3(new_n399), .A4(new_n372), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n371), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n394), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT77), .ZN(new_n404));
  OAI21_X1  g0204(.A(G169), .B1(new_n366), .B2(new_n367), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(KEYINPUT78), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI221_X1 g0208(.A(G169), .B1(KEYINPUT78), .B2(new_n406), .C1(new_n366), .C2(new_n367), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n368), .A2(G179), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n404), .A2(new_n400), .A3(new_n411), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n355), .A2(new_n402), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT82), .ZN(new_n414));
  INV_X1    g0214(.A(new_n271), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n256), .B2(G20), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n265), .A2(new_n416), .B1(new_n262), .B2(new_n415), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G58), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n373), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(new_n201), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT80), .ZN(new_n423));
  AOI21_X1  g0223(.A(G20), .B1(new_n341), .B2(new_n343), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(KEYINPUT7), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  OAI211_X1 g0226(.A(KEYINPUT80), .B(new_n426), .C1(new_n304), .C2(G20), .ZN(new_n427));
  AND2_X1   g0227(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n428));
  NOR2_X1   g0228(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n263), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n343), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n426), .A2(G20), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n425), .A2(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n422), .B1(new_n433), .B2(new_n373), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n270), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT79), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n342), .ZN(new_n438));
  NAND2_X1  g0238(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(G33), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n341), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n426), .A3(new_n221), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G68), .ZN(new_n443));
  AOI21_X1  g0243(.A(G20), .B1(new_n440), .B2(new_n341), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n426), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT16), .B(new_n422), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n418), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G87), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n228), .A2(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(G223), .B2(G1698), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n297), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n336), .A2(G232), .A3(new_n286), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n295), .A2(new_n453), .A3(KEYINPUT81), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n297), .A2(new_n300), .A3(new_n361), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n357), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n315), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n452), .A2(new_n457), .A3(new_n454), .A4(new_n369), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT17), .B1(new_n447), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n422), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n431), .A2(new_n432), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n342), .A2(G33), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n221), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT80), .B1(new_n467), .B2(new_n426), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n424), .A2(new_n423), .A3(KEYINPUT7), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n470), .B2(G68), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n264), .B(new_n446), .C1(new_n471), .C2(KEYINPUT16), .ZN(new_n472));
  AND4_X1   g0272(.A1(KEYINPUT17), .A2(new_n472), .A3(new_n417), .A4(new_n461), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n414), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n461), .A3(new_n417), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT17), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n447), .A2(KEYINPUT17), .A3(new_n461), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT82), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT18), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n458), .A2(G169), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n311), .B2(new_n458), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n447), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n472), .A2(new_n417), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT18), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n474), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n326), .A2(new_n413), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n440), .A2(new_n221), .A3(G68), .A4(new_n341), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT19), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n221), .B1(new_n360), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G87), .B2(new_n207), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n205), .B1(new_n272), .B2(new_n274), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n492), .B(new_n495), .C1(KEYINPUT19), .C2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n264), .B1(new_n262), .B2(new_n331), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n256), .A2(G33), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n261), .A2(new_n270), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n332), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G238), .A2(G1698), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n234), .B2(G1698), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n440), .A3(new_n341), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n336), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n299), .A2(G1), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n294), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G250), .B1(new_n299), .B2(G1), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n297), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n352), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n507), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n311), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n502), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(G190), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n261), .A2(new_n270), .A3(G87), .A4(new_n499), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n517), .B(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(G200), .B1(new_n507), .B2(new_n511), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n516), .A2(new_n519), .A3(new_n498), .A4(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n261), .A2(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n500), .B2(G97), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n276), .A2(G77), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT83), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n528), .A2(new_n205), .A3(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI221_X1 g0331(.A(new_n527), .B1(new_n221), .B2(new_n531), .C1(new_n433), .C2(new_n206), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n525), .B1(new_n532), .B2(new_n264), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n234), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n304), .A2(new_n305), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n304), .A2(G250), .A3(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n440), .A2(G244), .A3(new_n305), .A4(new_n341), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n534), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(KEYINPUT84), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n543), .A3(new_n534), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n336), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT85), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n298), .A3(KEYINPUT5), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT5), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(KEYINPUT85), .B2(G41), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n549), .A3(new_n508), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n356), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G257), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n336), .A2(new_n550), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(G200), .B1(new_n545), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n555), .ZN(new_n557));
  INV_X1    g0357(.A(new_n544), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n543), .B1(new_n540), .B2(new_n534), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n558), .A2(new_n559), .A3(new_n539), .ZN(new_n560));
  OAI211_X1 g0360(.A(G190), .B(new_n557), .C1(new_n560), .C2(new_n336), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n533), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n352), .B1(new_n545), .B2(new_n555), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n311), .B(new_n557), .C1(new_n560), .C2(new_n336), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n527), .B1(new_n221), .B2(new_n531), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n470), .B2(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n524), .B1(new_n566), .B2(new_n270), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n522), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G250), .A2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n553), .B2(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n440), .A3(new_n341), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n336), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n554), .A2(new_n235), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n311), .A3(new_n552), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n574), .A2(new_n575), .A3(new_n551), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(G169), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT23), .B1(new_n221), .B2(G107), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n206), .A3(G20), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n582), .C1(G20), .C2(new_n506), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT89), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  INV_X1    g0387(.A(G87), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n440), .A2(new_n221), .A3(new_n341), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n221), .A2(G87), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n344), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n585), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n264), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT25), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n261), .B2(G107), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n261), .A2(new_n598), .A3(G107), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT90), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(KEYINPUT90), .B(new_n598), .C1(new_n261), .C2(G107), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n500), .A2(G107), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n579), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n261), .A2(G116), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n500), .B2(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n229), .A2(G20), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n264), .A2(KEYINPUT88), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT88), .B1(new_n264), .B2(new_n611), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n538), .B(new_n221), .C1(G33), .C2(new_n205), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT20), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(KEYINPUT20), .B(new_n615), .C1(new_n612), .C2(new_n613), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n610), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n235), .A2(G1698), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G257), .B2(G1698), .ZN(new_n621));
  INV_X1    g0421(.A(G303), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n441), .A2(new_n621), .B1(new_n622), .B2(new_n304), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n551), .B1(new_n623), .B2(new_n297), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n554), .B2(new_n230), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n336), .A2(new_n550), .A3(KEYINPUT87), .A4(G270), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n352), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n619), .A2(KEYINPUT21), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n624), .A2(new_n628), .A3(G179), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT21), .B1(new_n619), .B2(new_n629), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n608), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n596), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n270), .B1(new_n636), .B2(new_n594), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n606), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n576), .A2(new_n552), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT91), .B1(new_n639), .B2(G190), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n578), .A2(new_n641), .A3(new_n369), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n640), .B(new_n642), .C1(G200), .C2(new_n578), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n624), .A2(new_n628), .A3(G190), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n624), .A2(new_n628), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n619), .B1(G200), .B2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n638), .A2(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n491), .A2(new_n569), .A3(new_n635), .A4(new_n647), .ZN(G372));
  AND3_X1   g0448(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT92), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT92), .B1(new_n484), .B2(new_n486), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n402), .A2(new_n474), .A3(new_n479), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n412), .A2(new_n354), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n323), .A2(new_n325), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n314), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n635), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n638), .A2(new_n643), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n569), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n515), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n515), .A2(new_n521), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n568), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n568), .B2(new_n664), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n491), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n659), .A2(new_n671), .ZN(G369));
  INV_X1    g0472(.A(new_n633), .ZN(new_n673));
  INV_X1    g0473(.A(new_n634), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n256), .A2(new_n221), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n619), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n675), .B(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n644), .B2(new_n646), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n681), .B1(new_n637), .B2(new_n606), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n608), .B1(new_n661), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n681), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n688), .B1(new_n608), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n608), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n675), .A2(new_n689), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n688), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(G399));
  NOR2_X1   g0496(.A1(new_n211), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n218), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n668), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n666), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n665), .A2(new_n703), .A3(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n663), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n662), .B1(new_n707), .B2(KEYINPUT94), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n568), .A2(new_n664), .A3(new_n667), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n703), .B2(new_n668), .ZN(new_n710));
  INV_X1    g0510(.A(new_n706), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n515), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT29), .B(new_n689), .C1(new_n708), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n670), .A2(new_n689), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n569), .A2(new_n635), .A3(new_n647), .A4(new_n689), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n576), .A2(new_n513), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n631), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n557), .B1(new_n560), .B2(new_n336), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n545), .A2(new_n555), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(KEYINPUT30), .A3(new_n631), .A4(new_n721), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n513), .A2(G179), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n723), .A2(new_n645), .A3(new_n639), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n681), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n719), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n715), .A2(new_n718), .B1(G330), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n702), .B1(new_n735), .B2(G1), .ZN(G364));
  INV_X1    g0536(.A(KEYINPUT96), .ZN(new_n737));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT95), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n256), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n737), .B1(new_n742), .B2(new_n697), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(KEYINPUT96), .A3(new_n698), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n211), .A2(new_n344), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G355), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G116), .B2(new_n210), .ZN(new_n749));
  INV_X1    g0549(.A(new_n441), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n211), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n299), .B2(new_n219), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n251), .A2(new_n299), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n220), .B1(G20), .B2(new_n352), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n746), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n221), .A2(new_n311), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n304), .B1(new_n765), .B2(new_n233), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n369), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n221), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n769), .A2(new_n202), .B1(new_n771), .B2(new_n588), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n315), .A2(G190), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n773), .A2(new_n221), .A3(new_n311), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n766), .B(new_n772), .C1(G58), .C2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(G20), .B1(new_n773), .B2(G179), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT98), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n770), .A2(new_n764), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n787));
  NAND3_X1  g0587(.A1(new_n770), .A2(new_n369), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n786), .A2(new_n787), .B1(G107), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n767), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n787), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G68), .A2(new_n791), .B1(new_n785), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n775), .A2(new_n782), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n780), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n774), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n798), .B1(new_n765), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n783), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n304), .B(new_n800), .C1(G329), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n771), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n768), .A2(G326), .B1(new_n803), .B2(G303), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n791), .A2(new_n805), .B1(new_n789), .B2(G283), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n794), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n762), .B1(new_n808), .B2(new_n759), .ZN(new_n809));
  INV_X1    g0609(.A(new_n758), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n684), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT99), .Z(new_n812));
  NOR2_X1   g0612(.A1(new_n686), .A2(new_n746), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G330), .B2(new_n684), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n335), .A2(new_n681), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n350), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n354), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n354), .A2(new_n681), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n716), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n817), .B2(new_n354), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n670), .A2(new_n689), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n734), .A2(G330), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n746), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n759), .A2(new_n756), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT100), .Z(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G77), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n797), .A2(new_n795), .B1(new_n783), .B2(new_n799), .ZN(new_n832));
  INV_X1    g0632(.A(new_n765), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n304), .B(new_n832), .C1(G116), .C2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n768), .A2(G303), .B1(new_n803), .B2(G107), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n788), .A2(new_n588), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G283), .B2(new_n791), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n782), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n788), .A2(new_n373), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n750), .B1(new_n840), .B2(new_n783), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G50), .C2(new_n803), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n833), .A2(G159), .B1(new_n774), .B2(G143), .ZN(new_n843));
  INV_X1    g0643(.A(new_n791), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n846), .C2(new_n769), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT34), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n842), .B(new_n849), .C1(new_n419), .C2(new_n780), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n847), .A2(new_n848), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n838), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n745), .B(new_n831), .C1(new_n852), .C2(new_n759), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n823), .B2(new_n757), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n828), .A2(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n740), .A2(new_n256), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT107), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT92), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n485), .A2(KEYINPUT18), .A3(new_n482), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT18), .B1(new_n485), .B2(new_n482), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n462), .A2(new_n473), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT92), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n447), .A2(new_n679), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n858), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n866), .ZN(new_n868));
  XOR2_X1   g0668(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n869));
  AND3_X1   g0669(.A1(new_n868), .A2(new_n475), .A3(new_n869), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n447), .A2(new_n483), .A3(KEYINPUT105), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n485), .B2(new_n482), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n859), .B1(new_n447), .B2(new_n483), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n485), .A2(KEYINPUT92), .A3(new_n482), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n868), .A2(new_n875), .A3(new_n475), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n869), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n870), .A2(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n865), .A2(new_n858), .A3(new_n866), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n445), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n373), .B1(new_n444), .B2(new_n426), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n463), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n264), .B1(new_n885), .B2(KEYINPUT16), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n886), .A2(KEYINPUT103), .B1(KEYINPUT16), .B2(new_n885), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n418), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n475), .B1(new_n889), .B2(new_n483), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n679), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n870), .A2(new_n874), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n488), .A2(KEYINPUT104), .A3(new_n891), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT104), .B1(new_n488), .B2(new_n891), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT38), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n857), .B1(new_n882), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n412), .A2(new_n681), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n824), .A2(new_n820), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n404), .A2(new_n400), .A3(new_n681), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n402), .A2(new_n412), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT102), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n404), .A2(new_n411), .A3(new_n400), .A4(new_n681), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n903), .A2(new_n897), .ZN(new_n915));
  INV_X1    g0715(.A(new_n651), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n914), .A2(new_n915), .B1(new_n916), .B2(new_n679), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n905), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n490), .B1(new_n717), .B2(new_n716), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n658), .B1(new_n715), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  INV_X1    g0721(.A(G330), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n911), .A2(new_n912), .ZN(new_n923));
  INV_X1    g0723(.A(new_n733), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT31), .B1(new_n729), .B2(new_n681), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n821), .B1(new_n926), .B2(new_n719), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT40), .B1(new_n915), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n865), .A2(new_n858), .A3(new_n866), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n931), .A2(new_n867), .A3(new_n879), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n897), .B1(new_n932), .B2(KEYINPUT38), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n927), .B(KEYINPUT40), .C1(new_n911), .C2(new_n912), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n930), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n490), .B1(new_n719), .B2(new_n926), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n922), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n856), .B1(new_n921), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n921), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n218), .A2(new_n233), .A3(new_n420), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n373), .A2(G50), .ZN(new_n943));
  OAI211_X1 g0743(.A(G1), .B(new_n738), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n531), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT35), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(G116), .A3(new_n222), .A4(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n944), .A3(new_n950), .ZN(G367));
  OAI211_X1 g0751(.A(new_n562), .B(new_n568), .C1(new_n533), .C2(new_n689), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n568), .B2(new_n689), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(KEYINPUT109), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(KEYINPUT109), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n957), .A2(new_n675), .A3(new_n689), .A4(new_n690), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT42), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n608), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n681), .B1(new_n960), .B2(new_n568), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT43), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n689), .B1(new_n519), .B2(new_n498), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n515), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n522), .B2(new_n964), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT108), .Z(new_n967));
  NAND3_X1  g0767(.A1(new_n962), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n963), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n963), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n959), .C2(new_n961), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n691), .A2(new_n956), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n697), .B(KEYINPUT41), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n956), .A2(new_n694), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n956), .A2(new_n694), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n977), .A2(new_n691), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n691), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n690), .B(new_n693), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n685), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n735), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n975), .B1(new_n989), .B2(new_n735), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n974), .B1(new_n990), .B2(new_n742), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n243), .A2(new_n752), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n760), .B1(new_n210), .B2(new_n331), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n746), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n844), .A2(new_n784), .B1(new_n419), .B2(new_n771), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n304), .B1(new_n783), .B2(new_n846), .C1(new_n202), .C2(new_n765), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n788), .A2(new_n233), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n781), .A2(G68), .ZN(new_n999));
  INV_X1    g0799(.A(G143), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(new_n1000), .B2(new_n769), .C1(new_n845), .C2(new_n797), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT111), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1002), .B2(new_n1001), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT112), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n844), .A2(new_n795), .B1(new_n788), .B2(new_n205), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n750), .B(new_n1006), .C1(G311), .C2(new_n768), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n803), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT46), .B1(new_n803), .B2(G116), .ZN(new_n1009));
  INV_X1    g0809(.A(G317), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n797), .A2(new_n622), .B1(new_n783), .B2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G283), .C2(new_n833), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n781), .A2(G107), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1008), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1005), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT47), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n994), .B1(new_n1016), .B2(new_n759), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n967), .A2(new_n758), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n991), .A2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n987), .A2(new_n988), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n697), .C1(new_n735), .C2(new_n985), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n699), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n747), .A2(new_n1023), .B1(new_n206), .B2(new_n211), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n247), .A2(new_n299), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n271), .A2(new_n202), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT50), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n699), .B(new_n299), .C1(new_n373), .C2(new_n233), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n751), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1024), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n745), .B1(new_n1030), .B2(new_n760), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n781), .A2(new_n332), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n202), .B2(new_n797), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT113), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n750), .B1(new_n373), .B2(new_n765), .C1(new_n845), .C2(new_n783), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n844), .A2(new_n415), .B1(new_n205), .B2(new_n788), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n769), .A2(new_n784), .B1(new_n771), .B2(new_n233), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n781), .A2(G283), .B1(G294), .B2(new_n803), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n833), .A2(G303), .B1(new_n774), .B2(G317), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n844), .B2(new_n799), .C1(new_n798), .C2(new_n769), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT114), .Z(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT115), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n750), .B1(G326), .B2(new_n801), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n229), .B2(new_n788), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1046), .B2(KEYINPUT49), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1038), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n759), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1031), .B1(new_n690), .B2(new_n810), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n985), .A2(new_n742), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1022), .A2(new_n1055), .ZN(G393));
  OAI21_X1  g0856(.A(new_n1021), .B1(new_n981), .B2(new_n982), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n697), .A3(new_n989), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n760), .B1(new_n205), .B2(new_n210), .C1(new_n752), .C2(new_n254), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n746), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n781), .A2(G77), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n769), .A2(new_n845), .B1(new_n784), .B2(new_n797), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n836), .B1(G50), .B2(new_n791), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n373), .B2(new_n771), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n415), .A2(new_n765), .B1(new_n1000), .B2(new_n783), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1067), .A2(new_n441), .A3(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n344), .B1(new_n783), .B2(new_n798), .C1(new_n795), .C2(new_n765), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n803), .A2(G283), .B1(new_n789), .B2(G107), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n622), .B2(new_n844), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G116), .C2(new_n781), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n768), .A2(G317), .B1(G311), .B2(new_n774), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n1065), .A2(new_n1069), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1060), .B1(new_n1052), .B2(new_n1076), .C1(new_n957), .C2(new_n810), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n983), .B2(new_n742), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1058), .A2(new_n1079), .ZN(G390));
  NAND3_X1  g0880(.A1(new_n734), .A2(G330), .A3(new_n823), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n908), .A2(new_n910), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT102), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n900), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n899), .A2(new_n904), .B1(new_n1086), .B2(new_n913), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n882), .B2(new_n898), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n689), .B(new_n818), .C1(new_n708), .C2(new_n714), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n923), .B1(new_n1089), .B2(new_n820), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1085), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n913), .A2(new_n1086), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n904), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n865), .A2(new_n866), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT107), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n879), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n881), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n902), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1099), .B2(new_n897), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1093), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n662), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n712), .B2(new_n713), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n707), .A2(KEYINPUT94), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n681), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n819), .B1(new_n1105), .B2(new_n818), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1086), .B(new_n933), .C1(new_n1106), .C2(new_n923), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n927), .B(G330), .C1(new_n911), .C2(new_n912), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1101), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1092), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1081), .A2(new_n1084), .A3(new_n1082), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1089), .A2(new_n820), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1081), .A2(new_n1084), .A3(new_n1082), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n906), .B1(new_n1113), .B2(new_n1085), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n490), .A2(new_n826), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1116), .B(new_n658), .C1(new_n715), .C2(new_n919), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT117), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT117), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1110), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1092), .A2(new_n1109), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1115), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1120), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n698), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n756), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n746), .B1(new_n271), .B2(new_n830), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n797), .A2(new_n229), .B1(new_n783), .B2(new_n795), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n304), .B(new_n1132), .C1(G97), .C2(new_n833), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n839), .B1(G87), .B2(new_n803), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G107), .A2(new_n791), .B1(new_n768), .B2(G283), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n1061), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n769), .A2(new_n1139), .B1(new_n788), .B2(new_n202), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G137), .B2(new_n791), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n803), .A2(G150), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n304), .B1(new_n797), .B2(new_n840), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n803), .B2(G150), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n765), .A2(new_n1146), .B1(new_n783), .B2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n781), .A2(G159), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1141), .A2(new_n1143), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1138), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1131), .B1(new_n1153), .B2(new_n759), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1130), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1124), .B2(new_n741), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1129), .A2(new_n1157), .ZN(G378));
  NOR2_X1   g0958(.A1(new_n285), .A2(new_n679), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n326), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n326), .A2(new_n1160), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n756), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n797), .A2(new_n206), .B1(new_n331), .B2(new_n765), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n750), .A2(G41), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G283), .C2(new_n801), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n788), .A2(new_n419), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G77), .B2(new_n803), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G97), .A2(new_n791), .B1(new_n768), .B2(G116), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n999), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G50), .B1(new_n263), .B2(new_n298), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1176), .A2(new_n1177), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n797), .A2(new_n1139), .B1(new_n765), .B2(new_n846), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G132), .B2(new_n791), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1146), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n768), .A2(G125), .B1(new_n803), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(new_n845), .C2(new_n780), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n789), .A2(G159), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n801), .C2(G124), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1179), .B1(new_n1177), .B2(new_n1176), .C1(new_n1185), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n759), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n745), .B1(new_n202), .B2(new_n829), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1168), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n935), .B1(new_n882), .B2(new_n898), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(G330), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1196), .A2(new_n930), .A3(new_n1167), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1167), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n488), .A2(new_n891), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT104), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n488), .A2(KEYINPUT104), .A3(new_n891), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT38), .B1(new_n1203), .B2(new_n894), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n929), .B1(new_n1204), .B2(new_n898), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT40), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n922), .B1(new_n933), .B2(new_n935), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1198), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n918), .B1(new_n1197), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1167), .B1(new_n1196), .B2(new_n930), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1198), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n905), .A4(new_n917), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1194), .B1(new_n1214), .B2(new_n742), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1117), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1197), .A2(new_n1209), .A3(new_n918), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1211), .A2(new_n1212), .B1(new_n905), .B2(new_n917), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n697), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1117), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1214), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1215), .B1(new_n1221), .B2(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n923), .A2(new_n756), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n750), .B1(new_n1139), .B2(new_n783), .C1(new_n845), .C2(new_n765), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1173), .B(new_n1226), .C1(G159), .C2(new_n803), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n791), .A2(new_n1182), .B1(G137), .B2(new_n774), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n840), .B2(new_n769), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT121), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1229), .A2(KEYINPUT121), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n781), .A2(G50), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1227), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n768), .A2(G294), .B1(new_n833), .B2(G107), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n229), .B2(new_n844), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT120), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n344), .B1(new_n783), .B2(new_n622), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G283), .B2(new_n774), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n997), .B1(G97), .B2(new_n803), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1032), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1052), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n830), .A2(G68), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1241), .A2(new_n745), .A3(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1115), .A2(new_n742), .B1(new_n1225), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n975), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1244), .B1(new_n1122), .B2(new_n1248), .ZN(G381));
  INV_X1    g1049(.A(G396), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1022), .A2(new_n1250), .A3(new_n1055), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1251), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G387), .A2(new_n1252), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n680), .A2(G213), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(G375), .A2(G378), .A3(new_n1254), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT122), .Z(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT124), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT60), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT60), .ZN(new_n1261));
  OAI211_X1 g1061(.A(KEYINPUT124), .B(new_n1261), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n697), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1245), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1246), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n698), .B1(new_n1259), .B2(KEYINPUT60), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(KEYINPUT125), .A4(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1244), .ZN(new_n1270));
  INV_X1    g1070(.A(G384), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(G384), .A3(new_n1244), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  INV_X1    g1074(.A(G2897), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1254), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1272), .A2(new_n1273), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1254), .A2(new_n1275), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1269), .B2(new_n1244), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1244), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1271), .B(new_n1281), .C1(new_n1265), .C2(new_n1268), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT123), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT123), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1210), .A2(new_n1213), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n742), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1222), .A2(new_n1247), .A3(new_n1214), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1193), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1156), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1215), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1254), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1251), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1250), .B1(new_n1022), .B2(new_n1055), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n991), .A2(G390), .A3(new_n1019), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G390), .B1(new_n991), .B2(new_n1019), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1303), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1299), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(KEYINPUT127), .A3(new_n1251), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1300), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1308), .A3(new_n1301), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1304), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1295), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1254), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(KEYINPUT63), .A3(new_n1312), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1296), .A2(new_n1310), .A3(new_n1314), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(new_n1316), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  AND4_X1   g1122(.A1(new_n1322), .A2(new_n1294), .A3(new_n1254), .A4(new_n1312), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1316), .B2(new_n1312), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1318), .B1(new_n1325), .B2(new_n1310), .ZN(G405));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1291), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1293), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1312), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1313), .A2(new_n1293), .A3(new_n1327), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1331), .A2(new_n1310), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1310), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


