//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT65), .B1(new_n461), .B2(new_n462), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n470), .A2(new_n476), .A3(G125), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n470), .A2(new_n476), .A3(KEYINPUT66), .A4(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n469), .B1(new_n482), .B2(G2105), .ZN(G160));
  NAND2_X1  g058(.A1(new_n464), .A2(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND2_X1   g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n465), .B(new_n492), .C1(new_n461), .C2(new_n462), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n470), .A2(new_n476), .A3(G138), .A4(new_n465), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT67), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n504), .A2(G543), .A3(new_n505), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n513), .A2(new_n502), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n511), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT68), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n504), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n507), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n520), .A2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(new_n509), .A2(G90), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n511), .A2(G52), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n502), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AOI22_X1  g109(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n502), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT69), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(G81), .B1(new_n511), .B2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT70), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G188));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT9), .B1(new_n518), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n511), .A2(new_n550), .A3(G53), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT71), .B(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n508), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n509), .A2(G91), .B1(G651), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G299));
  NAND2_X1  g132(.A1(G168), .A2(KEYINPUT72), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n559), .B1(new_n520), .B2(new_n527), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G286));
  OAI21_X1  g137(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n563));
  INV_X1    g138(.A(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n518), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n525), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n509), .A2(KEYINPUT73), .A3(G87), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n509), .A2(G86), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n511), .A2(G48), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n502), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n509), .A2(G85), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n511), .A2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n502), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n509), .A2(G92), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n508), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n511), .A2(G54), .B1(G651), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n582), .B1(new_n590), .B2(G868), .ZN(G284));
  OAI21_X1  g166(.A(new_n582), .B1(new_n590), .B2(G868), .ZN(G321));
  INV_X1    g167(.A(G299), .ZN(new_n593));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G286), .B2(new_n594), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT74), .ZN(G297));
  XOR2_X1   g172(.A(new_n596), .B(KEYINPUT75), .Z(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n539), .A2(new_n594), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n585), .A2(new_n589), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n603), .B2(new_n594), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g180(.A1(new_n470), .A2(new_n476), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n606), .A2(G2104), .A3(new_n465), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT13), .Z(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n464), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n486), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n465), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT78), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT77), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n631), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  AOI21_X1  g216(.A(KEYINPUT18), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2096), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G227));
  XOR2_X1   g222(.A(G1971), .B(G1976), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT19), .ZN(new_n649));
  XOR2_X1   g224(.A(G1956), .B(G2474), .Z(new_n650));
  XOR2_X1   g225(.A(G1961), .B(G1966), .Z(new_n651));
  AND2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n649), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n649), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G229));
  INV_X1    g239(.A(KEYINPUT36), .ZN(new_n665));
  INV_X1    g240(.A(G16), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G22), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(G166), .B2(new_n666), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT81), .B(G1971), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(G6), .A2(G16), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(G305), .B2(new_n666), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n666), .A2(G23), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n570), .B2(new_n666), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT33), .ZN(new_n679));
  INV_X1    g254(.A(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(new_n677), .C1(new_n570), .C2(new_n666), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n679), .B2(new_n682), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT83), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n676), .B(new_n687), .C1(new_n683), .C2(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n686), .A2(KEYINPUT34), .A3(new_n688), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G25), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n464), .A2(G131), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT79), .Z(new_n696));
  OAI21_X1  g271(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n697));
  INV_X1    g272(.A(G107), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G2105), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n486), .B2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n694), .B1(new_n702), .B2(new_n693), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT80), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n666), .A2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n666), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n691), .A2(new_n692), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n665), .B1(new_n712), .B2(KEYINPUT84), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n691), .A2(new_n714), .A3(new_n692), .A4(new_n711), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(KEYINPUT85), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n691), .A2(new_n665), .A3(new_n692), .A4(new_n711), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n713), .B2(new_n715), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n540), .A2(new_n666), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n666), .B2(G19), .ZN(new_n723));
  INV_X1    g298(.A(G1341), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n693), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n693), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT91), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n723), .A2(new_n724), .B1(G2090), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n666), .A2(G4), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n590), .B2(new_n666), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1348), .ZN(new_n733));
  INV_X1    g308(.A(G2078), .ZN(new_n734));
  NAND2_X1  g309(.A1(G164), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G27), .B2(G29), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n730), .B(new_n733), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G171), .A2(new_n666), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G5), .B2(new_n666), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT89), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n666), .A2(G21), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G168), .B2(new_n666), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n666), .A2(G20), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT23), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  INV_X1    g326(.A(G1956), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(G160), .A2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G34), .Z(new_n756));
  OAI21_X1  g331(.A(new_n754), .B1(G29), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n723), .A2(new_n724), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n606), .A2(G127), .ZN(new_n762));
  NAND2_X1  g337(.A1(G115), .A2(G2104), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n465), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT86), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  AOI211_X1 g342(.A(new_n764), .B(new_n767), .C1(G139), .C2(new_n464), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n693), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n693), .B2(G33), .ZN(new_n770));
  INV_X1    g345(.A(G2072), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n770), .A2(new_n771), .B1(new_n740), .B2(new_n739), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n693), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n464), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n486), .A2(G128), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n693), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n784), .A2(new_n693), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n617), .B2(new_n693), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n693), .A2(G32), .ZN(new_n790));
  NAND3_X1  g365(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT88), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT26), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n486), .A2(G129), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n693), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT27), .B(G1996), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n729), .A2(G2090), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n736), .A2(new_n734), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n789), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AND4_X1   g377(.A1(new_n761), .A2(new_n772), .A3(new_n773), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n737), .A2(new_n748), .A3(new_n760), .A4(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n717), .A2(new_n721), .A3(new_n804), .ZN(G311));
  NOR2_X1   g380(.A1(new_n721), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n716), .ZN(G150));
  NAND2_X1  g382(.A1(new_n511), .A2(G55), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT92), .B(G93), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(new_n502), .B2(new_n809), .C1(new_n525), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G860), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n590), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n811), .B(new_n539), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G860), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n821), .B(new_n822), .C1(new_n818), .C2(new_n817), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n819), .A2(new_n820), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n813), .B1(new_n823), .B2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n781), .B(G164), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n768), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n796), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n701), .B(new_n608), .ZN(new_n830));
  OR2_X1    g405(.A1(G106), .A2(G2105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n832));
  INV_X1    g407(.A(G130), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n485), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G142), .B2(new_n464), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n828), .A2(new_n829), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(G160), .B(new_n617), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G162), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n828), .B(new_n836), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n839), .C1(new_n840), .C2(new_n829), .ZN(new_n841));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n841), .B(new_n842), .C1(new_n840), .C2(new_n839), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g419(.A1(new_n811), .A2(new_n594), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n570), .A2(new_n708), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n570), .A2(new_n708), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(KEYINPUT95), .A3(new_n847), .ZN(new_n852));
  XNOR2_X1  g427(.A(G303), .B(G305), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(new_n846), .C1(new_n849), .C2(new_n848), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT42), .ZN(new_n858));
  INV_X1    g433(.A(new_n816), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n603), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n590), .A2(new_n593), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n602), .A2(G299), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n861), .B2(new_n862), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n864), .B1(new_n868), .B2(new_n860), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n858), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n845), .B1(new_n870), .B2(new_n594), .ZN(G295));
  OAI21_X1  g446(.A(new_n845), .B1(new_n870), .B2(new_n594), .ZN(G331));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n561), .A2(G171), .ZN(new_n874));
  INV_X1    g449(.A(G168), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G301), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n859), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  AOI21_X1  g453(.A(G301), .B1(new_n558), .B2(new_n560), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n816), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n859), .A2(new_n874), .A3(KEYINPUT97), .A4(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n863), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n887), .B(new_n816), .C1(new_n878), .C2(new_n879), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n877), .A2(new_n880), .A3(KEYINPUT96), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n868), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n857), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n842), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n854), .A2(new_n856), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n854), .B2(new_n856), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n863), .B(new_n865), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n863), .B1(new_n889), .B2(new_n888), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT100), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n897), .B(new_n903), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n893), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n873), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n893), .ZN(new_n908));
  INV_X1    g483(.A(new_n904), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n889), .A2(new_n888), .ZN(new_n910));
  OAI22_X1  g485(.A1(new_n910), .A2(new_n863), .B1(new_n898), .B2(new_n884), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n903), .B1(new_n911), .B2(new_n897), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n908), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n895), .A2(new_n896), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n886), .A2(new_n890), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(KEYINPUT98), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT98), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n886), .A2(new_n890), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n893), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n915), .B1(new_n921), .B2(new_n906), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n907), .A2(new_n914), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n908), .B(new_n906), .C1(new_n909), .C2(new_n912), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n921), .B2(new_n906), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n915), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(G397));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(G160), .B2(G40), .ZN(new_n928));
  INV_X1    g503(.A(new_n481), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n477), .B2(new_n478), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n465), .B1(new_n930), .B2(new_n480), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n932));
  INV_X1    g507(.A(G40), .ZN(new_n933));
  NOR4_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n469), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G164), .B2(G1384), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n928), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G1986), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n708), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT103), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n938), .B2(new_n708), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n701), .B(new_n704), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(KEYINPUT104), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n796), .B(G1996), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n780), .B(G2067), .Z(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(KEYINPUT104), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n937), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n500), .A2(new_n499), .ZN(new_n952));
  INV_X1    g527(.A(new_n498), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR4_X1   g531(.A1(G164), .A2(KEYINPUT105), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n482), .A2(G2105), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G40), .A3(new_n468), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n932), .ZN(new_n961));
  NAND3_X1  g536(.A1(G160), .A2(KEYINPUT102), .A3(G40), .ZN(new_n962));
  INV_X1    g537(.A(new_n954), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n958), .A2(new_n961), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT115), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n928), .A2(new_n934), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n964), .A4(new_n958), .ZN(new_n969));
  INV_X1    g544(.A(G1348), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n961), .A2(new_n954), .A3(new_n962), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(G2067), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT60), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n590), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n590), .A2(new_n975), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n978), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n971), .A2(new_n973), .A3(new_n980), .A4(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n971), .A2(new_n973), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n974), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n988));
  NOR3_X1   g563(.A1(G164), .A2(new_n935), .A3(G1384), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT56), .B(G2072), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n967), .A2(new_n987), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n954), .A2(new_n955), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n961), .A2(new_n962), .A3(new_n964), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n752), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n961), .A2(new_n962), .A3(new_n990), .A4(new_n991), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT113), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n552), .A2(new_n998), .A3(new_n556), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n552), .B2(new_n556), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n992), .A2(new_n995), .A3(new_n997), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(KEYINPUT113), .A2(new_n996), .B1(new_n994), .B2(new_n752), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(KEYINPUT114), .A3(new_n1001), .A4(new_n992), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n992), .A2(new_n995), .A3(new_n997), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1001), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n979), .A2(new_n983), .A3(KEYINPUT118), .A4(new_n981), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(KEYINPUT61), .A3(new_n1002), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n936), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n928), .A2(new_n934), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT58), .B(G1341), .Z(new_n1021));
  AOI22_X1  g596(.A1(new_n1019), .A2(new_n1020), .B1(new_n972), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1022), .B2(new_n539), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n972), .A2(new_n1021), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n961), .A2(new_n962), .A3(new_n990), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G1996), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT116), .B(new_n540), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1027), .A3(KEYINPUT59), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1016), .B(new_n1029), .C1(new_n1022), .C2(new_n539), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1015), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n986), .A2(new_n1013), .A3(new_n1014), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n982), .A2(new_n590), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1010), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1007), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1018), .A2(new_n1037), .A3(G2078), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n960), .A2(KEYINPUT122), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n960), .A2(KEYINPUT122), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT123), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n966), .A2(new_n969), .A3(new_n740), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1025), .B2(G2078), .ZN(new_n1045));
  XOR2_X1   g620(.A(G301), .B(KEYINPUT54), .Z(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n967), .A2(new_n1038), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1046), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n967), .A2(new_n758), .A3(new_n964), .A4(new_n958), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1025), .A2(new_n745), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G168), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1053), .A2(new_n1061), .A3(new_n1054), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n875), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1066), .A2(KEYINPUT120), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(KEYINPUT120), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1060), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1052), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n1073));
  OAI22_X1  g648(.A1(G166), .A2(new_n1057), .B1(KEYINPUT106), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT106), .B(KEYINPUT55), .Z(new_n1075));
  NAND3_X1  g650(.A1(G303), .A2(G8), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n965), .A2(G2090), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1019), .A2(G1971), .ZN(new_n1079));
  OAI211_X1 g654(.A(G8), .B(new_n1077), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1079), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n994), .A2(G2090), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1057), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1083), .B2(new_n1077), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(new_n680), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n680), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT107), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n972), .A2(new_n1088), .A3(G8), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n972), .B2(G8), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1086), .B(new_n1087), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G305), .A2(G1981), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n572), .A2(new_n573), .A3(new_n1093), .A4(new_n575), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT49), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n928), .A2(new_n934), .A3(new_n963), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT107), .B1(new_n1098), .B2(new_n1057), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n972), .A2(new_n1088), .A3(G8), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1085), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1091), .B(new_n1097), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT109), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT52), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1107), .A2(KEYINPUT109), .A3(new_n1091), .A4(new_n1097), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1084), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1072), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1036), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1055), .A2(KEYINPUT119), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(G168), .A3(new_n1062), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1069), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1114), .A2(new_n1115), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1071), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1112), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1049), .A2(G171), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1084), .B(new_n1121), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1097), .A2(new_n680), .A3(new_n570), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1126), .A2(new_n1094), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT108), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1103), .B(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1080), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1111), .A2(new_n1125), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1055), .A2(G8), .A3(new_n561), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1084), .B(new_n1133), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT110), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT63), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1109), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT110), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1137), .A2(KEYINPUT63), .ZN(new_n1140));
  OAI21_X1  g715(.A(G8), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1074), .A2(KEYINPUT111), .A3(new_n1076), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1103), .A2(new_n1128), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1103), .A2(new_n1128), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1140), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT112), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1129), .A2(KEYINPUT112), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1136), .A2(new_n1139), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n950), .B1(new_n1132), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n937), .A2(new_n1020), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT46), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n946), .A2(new_n796), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1152), .A2(new_n1153), .B1(new_n937), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT47), .ZN(new_n1157));
  INV_X1    g732(.A(new_n937), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n780), .A2(G2067), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n702), .A2(new_n704), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT125), .Z(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1161), .B2(new_n947), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT48), .B1(new_n940), .B2(new_n937), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n940), .A2(KEYINPUT48), .A3(new_n937), .ZN(new_n1164));
  INV_X1    g739(.A(new_n949), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1158), .ZN(new_n1166));
  OAI221_X1 g741(.A(new_n1157), .B1(new_n1158), .B2(new_n1162), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT126), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1151), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g744(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1171));
  XNOR2_X1  g745(.A(new_n1171), .B(KEYINPUT127), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n1172), .A3(new_n843), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


