//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n201), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n219), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n214), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  AND2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G1698), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G222), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n251), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n256), .A3(G274), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(KEYINPUT65), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT65), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n264), .A2(new_n256), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n263), .B1(new_n269), .B2(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n258), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n226), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n226), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT66), .B1(G20), .B2(G33), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n274), .B1(new_n275), .B2(new_n276), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n225), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n226), .A3(G1), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n285), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n208), .B1(new_n265), .B2(G20), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(new_n290), .B1(new_n208), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n258), .A2(new_n293), .A3(new_n270), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n273), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n271), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n258), .A2(G190), .A3(new_n270), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n286), .A2(KEYINPUT9), .A3(new_n291), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n297), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n299), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n300), .A4(new_n297), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n249), .A2(G232), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n309));
  INV_X1    g0109(.A(G107), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n251), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n257), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n263), .B1(new_n269), .B2(G244), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n272), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n281), .A2(new_n275), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n317), .A2(new_n276), .B1(new_n226), .B2(new_n253), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n285), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n253), .B1(new_n265), .B2(G20), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n289), .A2(new_n320), .B1(new_n253), .B2(new_n288), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n315), .B(new_n322), .C1(G179), .C2(new_n314), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n314), .A2(G200), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n312), .A2(G190), .A3(new_n313), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n319), .A3(new_n321), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n296), .A2(new_n307), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  OR2_X1    g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n226), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n332), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n202), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G58), .A2(G68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT71), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(G58), .A3(G68), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(new_n203), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G20), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n279), .A2(new_n280), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G159), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n330), .B1(new_n337), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n202), .B1(new_n333), .B2(KEYINPUT7), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n246), .A2(new_n247), .A3(G20), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n334), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(G20), .A2(new_n342), .B1(new_n344), .B2(G159), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n285), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n275), .B1(new_n265), .B2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n289), .B1(new_n288), .B2(new_n275), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT18), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n264), .A2(G232), .A3(new_n268), .A4(new_n256), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G223), .A2(G1698), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n209), .B2(G1698), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n251), .B1(G33), .B2(G87), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n359), .B(new_n262), .C1(new_n362), .C2(new_n256), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G169), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n293), .B2(new_n363), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n357), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n358), .B1(new_n357), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT72), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n363), .A2(G200), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n354), .A2(new_n370), .A3(new_n356), .A4(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(new_n365), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n358), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n368), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n226), .A2(G68), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n380), .B1(new_n253), .B2(new_n276), .C1(new_n281), .C2(new_n208), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT68), .B1(new_n381), .B2(new_n285), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT11), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n281), .A2(new_n208), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n380), .B1(new_n276), .B2(new_n253), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT68), .B(new_n285), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n387), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT11), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n287), .A2(G1), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT12), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n379), .C1(KEYINPUT69), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(KEYINPUT69), .ZN(new_n394));
  XOR2_X1   g0194(.A(new_n393), .B(new_n394), .Z(new_n395));
  AOI21_X1  g0195(.A(new_n202), .B1(new_n265), .B2(G20), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n289), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n388), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n214), .A2(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G226), .B2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n401), .B2(new_n248), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n263), .B1(new_n402), .B2(new_n257), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n269), .A2(G238), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n403), .B2(new_n404), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n407), .A2(new_n369), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G200), .ZN(new_n410));
  INV_X1    g0210(.A(new_n408), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(new_n406), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n398), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n407), .A2(new_n408), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT14), .B1(new_n414), .B2(new_n272), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(G179), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n406), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(G169), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n413), .B1(new_n420), .B2(new_n398), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n329), .A2(new_n378), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n260), .A2(G1), .ZN(new_n424));
  AND2_X1   g0224(.A1(KEYINPUT5), .A2(G41), .ZN(new_n425));
  NOR2_X1   g0225(.A1(KEYINPUT5), .A2(G41), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(G264), .A3(new_n256), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT5), .B(G41), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(G274), .A3(new_n256), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(G257), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n433));
  INV_X1    g0233(.A(G1698), .ZN(new_n434));
  OAI211_X1 g0234(.A(G250), .B(new_n434), .C1(new_n246), .C2(new_n247), .ZN(new_n435));
  INV_X1    g0235(.A(G294), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n433), .B(new_n435), .C1(new_n278), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT82), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n437), .A2(new_n438), .A3(new_n257), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n437), .B2(new_n257), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n369), .B(new_n432), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n257), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n410), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT79), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n226), .B(G87), .C1(new_n246), .C2(new_n247), .ZN(new_n447));
  AND2_X1   g0247(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n446), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(G20), .B1(new_n331), .B2(new_n332), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n448), .A2(new_n449), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(KEYINPUT79), .A3(G87), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n447), .A2(KEYINPUT22), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT24), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT23), .B1(new_n226), .B2(G107), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n310), .A3(G20), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n456), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n457), .B1(new_n456), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n285), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n391), .A2(G20), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT25), .ZN(new_n469));
  AOI211_X1 g0269(.A(G107), .B(new_n468), .C1(KEYINPUT81), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(KEYINPUT81), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n278), .A2(G1), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n288), .A2(new_n285), .A3(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n472), .A2(new_n473), .B1(G107), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n445), .A2(new_n467), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G169), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n431), .B1(new_n257), .B2(new_n437), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G179), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n467), .A2(new_n476), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT74), .ZN(new_n484));
  INV_X1    g0284(.A(new_n285), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT6), .ZN(new_n486));
  AND2_X1   g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G97), .A2(G107), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT6), .A2(G97), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT73), .B1(new_n490), .B2(G107), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT73), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n310), .A3(KEYINPUT6), .A4(G97), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(G20), .B1(G77), .B2(new_n344), .ZN(new_n495));
  XOR2_X1   g0295(.A(KEYINPUT70), .B(KEYINPUT7), .Z(new_n496));
  OAI21_X1  g0296(.A(new_n336), .B1(new_n349), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G107), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n485), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n468), .A2(G97), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n475), .B2(G97), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n484), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n494), .A2(G20), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n344), .A2(G77), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n310), .B1(new_n335), .B2(new_n336), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n285), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n501), .A3(KEYINPUT74), .ZN(new_n509));
  OAI211_X1 g0309(.A(G244), .B(new_n434), .C1(new_n246), .C2(new_n247), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n434), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n512), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n257), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n427), .A2(new_n256), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n216), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AND4_X1   g0320(.A1(new_n369), .A2(new_n517), .A3(new_n430), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n516), .B2(new_n257), .ZN(new_n522));
  AOI21_X1  g0322(.A(G200), .B1(new_n522), .B2(new_n430), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n503), .B(new_n509), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n522), .A2(G179), .A3(new_n430), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n272), .B1(new_n522), .B2(new_n430), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(new_n499), .B2(new_n502), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(G264), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(new_n434), .C1(new_n246), .C2(new_n247), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n331), .A2(G303), .A3(new_n332), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n257), .ZN(new_n533));
  INV_X1    g0333(.A(new_n225), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n429), .A2(new_n424), .B1(new_n534), .B2(new_n255), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT77), .B1(new_n535), .B2(G270), .ZN(new_n536));
  AND4_X1   g0336(.A1(KEYINPUT77), .A2(new_n427), .A3(G270), .A4(new_n256), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n430), .B(new_n533), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  INV_X1    g0339(.A(new_n430), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT77), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n518), .B2(new_n211), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n535), .A2(KEYINPUT77), .A3(G270), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(G190), .A3(new_n533), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n514), .B(new_n226), .C1(G33), .C2(new_n215), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n210), .A2(G20), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n285), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT20), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n546), .A2(KEYINPUT20), .A3(new_n285), .A4(new_n547), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n468), .A2(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n475), .B2(G116), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n539), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n272), .B1(new_n552), .B2(new_n554), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n538), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n538), .A2(new_n558), .A3(KEYINPUT21), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n544), .A2(new_n555), .A3(G179), .A4(new_n533), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n226), .B1(new_n399), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n488), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n452), .A2(G68), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT76), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n566), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n565), .B1(new_n276), .B2(new_n215), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n570), .A2(new_n571), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n285), .B1(new_n288), .B2(new_n317), .ZN(new_n576));
  INV_X1    g0376(.A(new_n317), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n475), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT75), .ZN(new_n580));
  OR2_X1    g0380(.A1(G238), .A2(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(G244), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G1698), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n583), .C1(new_n246), .C2(new_n247), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G116), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n257), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n256), .A2(G274), .A3(new_n424), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n265), .A2(G45), .ZN(new_n589));
  AND2_X1   g0389(.A1(G33), .A2(G41), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(G250), .C1(new_n590), .C2(new_n225), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G169), .B1(new_n587), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n256), .B1(new_n584), .B2(new_n585), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n592), .A3(G179), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n580), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n587), .A2(new_n593), .A3(new_n293), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n595), .A2(new_n592), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(KEYINPUT75), .C1(G169), .C2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n579), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n599), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n475), .A2(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(G190), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n576), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n564), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n423), .A2(new_n483), .A3(new_n528), .A4(new_n608), .ZN(new_n609));
  XOR2_X1   g0409(.A(new_n609), .B(KEYINPUT83), .Z(G372));
  INV_X1    g0410(.A(new_n367), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n357), .A2(new_n358), .A3(new_n365), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n420), .A2(new_n398), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n413), .B2(new_n323), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n373), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n307), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT87), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n592), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n588), .A2(KEYINPUT84), .A3(new_n591), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n595), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(KEYINPUT85), .B(new_n598), .C1(new_n625), .C2(G169), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n588), .A2(KEYINPUT84), .A3(new_n591), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT84), .B1(new_n588), .B2(new_n591), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n587), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n272), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT85), .B1(new_n631), .B2(new_n598), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n579), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n482), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n445), .A2(new_n467), .A3(new_n476), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(G200), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n576), .A3(new_n604), .A4(new_n605), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n524), .A3(new_n527), .A4(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n633), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n607), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT86), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n517), .A2(new_n430), .A3(new_n520), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G169), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n522), .A2(G179), .A3(new_n430), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n508), .B2(new_n501), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT26), .A4(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n503), .A2(new_n509), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n633), .A3(new_n638), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n646), .A2(KEYINPUT26), .A3(new_n606), .A4(new_n601), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n649), .A2(new_n650), .B1(new_n651), .B2(KEYINPUT86), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n640), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  OAI221_X1 g0453(.A(new_n296), .B1(new_n616), .B2(new_n621), .C1(new_n422), .C2(new_n653), .ZN(G369));
  NAND2_X1  g0454(.A1(new_n391), .A2(new_n226), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n555), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n634), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n663), .B(KEYINPUT88), .C1(new_n564), .C2(new_n662), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(KEYINPUT88), .B2(new_n663), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT89), .Z(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n467), .ZN(new_n668));
  INV_X1    g0468(.A(new_n476), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n660), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n483), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n479), .A2(new_n481), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n668), .B2(new_n669), .ZN(new_n673));
  INV_X1    g0473(.A(new_n660), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n634), .A2(new_n674), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT90), .Z(new_n678));
  AND2_X1   g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n482), .B2(new_n674), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n222), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  NOR4_X1   g0483(.A1(new_n683), .A2(new_n265), .A3(G116), .A4(new_n568), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n229), .B2(new_n683), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT28), .Z(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n653), .B2(new_n660), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n649), .A2(new_n650), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n651), .A2(KEYINPUT86), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n647), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n633), .ZN(new_n693));
  AND4_X1   g0493(.A1(new_n636), .A2(new_n524), .A3(new_n527), .A4(new_n638), .ZN(new_n694));
  INV_X1    g0494(.A(new_n634), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n673), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT94), .A3(new_n674), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n688), .A2(new_n689), .A3(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n607), .A2(new_n527), .A3(KEYINPUT26), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(KEYINPUT26), .B2(new_n649), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n660), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(new_n689), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g0505(.A(KEYINPUT92), .B(KEYINPUT30), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n538), .A2(new_n293), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n443), .A2(new_n602), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .A4(new_n522), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n522), .A2(new_n480), .A3(new_n599), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n544), .A2(G179), .A3(new_n533), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT91), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n706), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n707), .A2(new_n522), .A3(new_n709), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(new_n643), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT93), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n630), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n432), .B2(new_n442), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n587), .B(KEYINPUT93), .C1(new_n628), .C2(new_n629), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n538), .A4(new_n721), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n660), .B1(new_n714), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n483), .A2(new_n608), .A3(new_n528), .A4(new_n674), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT31), .B(new_n660), .C1(new_n714), .C2(new_n723), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n705), .B1(G330), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n686), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n287), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n265), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n683), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n667), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n666), .ZN(new_n737));
  INV_X1    g0537(.A(new_n735), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n225), .B1(G20), .B2(new_n272), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n222), .A2(G355), .A3(new_n251), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G116), .B2(new_n222), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n682), .A2(new_n251), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n260), .B2(new_n229), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n241), .A2(new_n260), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n742), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n226), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n369), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n248), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n369), .A2(new_n410), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n757), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n226), .A2(new_n293), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G303), .A2(new_n763), .B1(new_n767), .B2(G311), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n764), .A2(new_n761), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n226), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n760), .B(new_n771), .C1(G294), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n764), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n776), .A2(new_n410), .A3(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT33), .B(G317), .Z(new_n779));
  NOR3_X1   g0579(.A1(new_n776), .A2(new_n369), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n778), .A2(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n757), .A2(new_n765), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G329), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n775), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n758), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G107), .A2(new_n792), .B1(new_n763), .B2(G87), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n253), .B2(new_n766), .C1(new_n201), .C2(new_n781), .ZN(new_n794));
  INV_X1    g0594(.A(new_n770), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n248), .B(new_n794), .C1(G50), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OR3_X1    g0597(.A1(new_n788), .A2(KEYINPUT32), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(KEYINPUT32), .B1(new_n788), .B2(new_n797), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G68), .A2(new_n777), .B1(new_n774), .B2(G97), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT97), .Z(new_n802));
  OAI21_X1  g0602(.A(new_n791), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n756), .B1(new_n803), .B2(new_n746), .ZN(new_n804));
  INV_X1    g0604(.A(new_n745), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n666), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n737), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n323), .A2(new_n660), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n322), .A2(new_n660), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n326), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n323), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n688), .B2(new_n699), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n328), .A2(new_n674), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n692), .B2(new_n697), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n729), .A2(G330), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n735), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n746), .A2(new_n743), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n741), .B1(new_n253), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n746), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n248), .B1(new_n758), .B2(new_n567), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G303), .A2(new_n795), .B1(new_n767), .B2(G116), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n310), .B2(new_n762), .C1(new_n759), .C2(new_n778), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(G311), .C2(new_n789), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G294), .A2(new_n780), .B1(new_n774), .B2(G97), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT99), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n777), .A2(G150), .B1(new_n795), .B2(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n781), .C1(new_n797), .C2(new_n766), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT34), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G68), .A2(new_n792), .B1(new_n763), .B2(G50), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n788), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n251), .B1(new_n773), .B2(new_n201), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n826), .A2(new_n828), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n821), .B1(new_n822), .B2(new_n840), .C1(new_n812), .C2(new_n744), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n819), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  OR2_X1    g0643(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n844), .A2(G116), .A3(new_n227), .A4(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT36), .Z(new_n847));
  NAND4_X1  g0647(.A1(new_n229), .A2(G77), .A3(new_n341), .A4(new_n339), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n208), .A2(G68), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n265), .B(G13), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n658), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT102), .B1(new_n357), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT102), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n854), .B(new_n658), .C1(new_n354), .C2(new_n356), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n374), .B(new_n372), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n357), .A2(new_n852), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n357), .A2(KEYINPUT102), .A3(new_n852), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n374), .A2(new_n372), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n370), .A2(new_n371), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n865), .A2(KEYINPUT17), .A3(new_n354), .A4(new_n356), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT17), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n372), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n613), .A2(new_n869), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n857), .A2(new_n864), .B1(new_n870), .B2(new_n862), .ZN(new_n871));
  XNOR2_X1  g0671(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n353), .A2(new_n285), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT16), .B1(new_n351), .B2(new_n352), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n356), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n365), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n852), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n372), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n882));
  INV_X1    g0682(.A(new_n878), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n377), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT103), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n880), .C1(new_n856), .C2(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT38), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n873), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n882), .A2(new_n886), .A3(new_n884), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n420), .A2(new_n398), .A3(new_n674), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n890), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n413), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n398), .A2(new_n660), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n614), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n398), .B(new_n660), .C1(new_n413), .C2(new_n420), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n815), .B2(new_n809), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT101), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT101), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n902), .C1(new_n815), .C2(new_n809), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n893), .A2(new_n887), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n613), .A2(new_n658), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n897), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n422), .B1(new_n700), .B2(new_n704), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n296), .B1(new_n616), .B2(new_n621), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n910), .B(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  AND4_X1   g0715(.A1(new_n915), .A2(new_n729), .A3(new_n902), .A4(new_n812), .ZN(new_n916));
  INV_X1    g0716(.A(new_n887), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n881), .A2(KEYINPUT103), .B1(new_n377), .B2(new_n883), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n918), .B2(new_n886), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n729), .A2(new_n902), .A3(new_n812), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n887), .B2(new_n873), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n423), .A3(new_n729), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n729), .A2(new_n902), .A3(new_n812), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n915), .B1(new_n888), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n729), .A2(new_n902), .A3(new_n812), .A4(new_n915), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n893), .B2(new_n887), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n423), .A2(new_n729), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(G330), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n914), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n265), .B2(new_n732), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n914), .A2(new_n932), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n851), .B1(new_n934), .B2(new_n935), .ZN(G367));
  AND2_X1   g0736(.A1(new_n751), .A2(new_n237), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n747), .B1(new_n222), .B2(new_n317), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n758), .A2(new_n215), .ZN(new_n939));
  INV_X1    g0739(.A(G303), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n436), .A2(new_n778), .B1(new_n781), .B2(new_n940), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(G311), .C2(new_n795), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n762), .A2(new_n210), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n251), .B(new_n944), .C1(G283), .C2(new_n767), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G107), .A2(new_n774), .B1(new_n943), .B2(KEYINPUT46), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n789), .A2(G317), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n942), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n780), .A2(G150), .B1(G50), .B2(new_n767), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n792), .A2(G77), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n949), .A2(new_n251), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n773), .A2(new_n202), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n789), .A2(G137), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n770), .A2(new_n830), .B1(new_n762), .B2(new_n201), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G159), .B2(new_n777), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n951), .A2(new_n953), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT47), .Z(new_n959));
  OAI221_X1 g0759(.A(new_n742), .B1(new_n937), .B2(new_n938), .C1(new_n959), .C2(new_n822), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT111), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n633), .A2(new_n638), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n576), .A2(new_n604), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n660), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n693), .B2(new_n964), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT105), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n745), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n503), .A2(new_n509), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n528), .B1(new_n970), .B2(new_n674), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n648), .A2(new_n660), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n680), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n680), .A2(new_n973), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n676), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n667), .B(new_n675), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n678), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n730), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(new_n730), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n683), .B(KEYINPUT41), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n733), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n967), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT108), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n967), .A2(new_n987), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n989), .B1(KEYINPUT109), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n679), .A2(new_n973), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT107), .ZN(new_n995));
  INV_X1    g0795(.A(new_n973), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n527), .B1(new_n996), .B2(new_n673), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n993), .A2(KEYINPUT42), .B1(new_n674), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT106), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n992), .A2(new_n1002), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n1003), .A2(new_n676), .A3(new_n996), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n676), .B2(new_n996), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n969), .B1(new_n986), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(G387));
  OR2_X1    g0810(.A1(new_n982), .A2(new_n730), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n982), .A2(new_n730), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n683), .A3(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n675), .A2(new_n805), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n234), .A2(G45), .A3(new_n248), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT50), .B1(new_n275), .B2(G50), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1016), .B(new_n260), .C1(new_n202), .C2(new_n253), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n275), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n248), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1019), .A2(new_n567), .A3(new_n210), .A4(new_n488), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n682), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n747), .B1(new_n222), .B2(new_n310), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n742), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n773), .A2(new_n317), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G50), .B2(new_n780), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT112), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n778), .A2(new_n275), .B1(new_n770), .B2(new_n797), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n202), .A2(new_n766), .B1(new_n762), .B2(new_n253), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n248), .A4(new_n939), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1026), .B(new_n1029), .C1(new_n282), .C2(new_n788), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n774), .A2(G283), .B1(new_n763), .B2(G294), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n780), .A2(G317), .B1(G303), .B2(new_n767), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n777), .A2(G311), .B1(new_n795), .B2(G322), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT113), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT49), .Z(new_n1040));
  OAI221_X1 g0840(.A(new_n248), .B1(new_n210), .B2(new_n758), .C1(new_n788), .C2(new_n769), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1023), .B1(new_n1042), .B2(new_n746), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n982), .A2(new_n734), .B1(new_n1014), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1013), .A2(new_n1044), .ZN(G393));
  INV_X1    g0845(.A(new_n980), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n1012), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(new_n683), .A3(new_n983), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n996), .A2(new_n745), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n752), .A2(new_n244), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n747), .B1(new_n222), .B2(new_n215), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n742), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n780), .A2(G159), .B1(new_n795), .B2(G150), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n763), .A2(G68), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n275), .B2(new_n766), .C1(new_n778), .C2(new_n208), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n773), .A2(new_n253), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n251), .C1(new_n567), .C2(new_n758), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1054), .B(new_n1060), .C1(new_n830), .C2(new_n788), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n780), .A2(G311), .B1(new_n795), .B2(G317), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  AOI22_X1  g0863(.A1(G303), .A2(new_n777), .B1(new_n774), .B2(G116), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT115), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(new_n436), .C2(new_n766), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n251), .B1(new_n792), .B2(G107), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n759), .B2(new_n762), .C1(new_n788), .C2(new_n782), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT114), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1061), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1052), .B1(new_n1070), .B2(new_n746), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n980), .A2(new_n734), .B1(new_n1049), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1048), .A2(new_n1072), .ZN(G390));
  NOR2_X1   g0873(.A1(new_n817), .A2(new_n422), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n911), .A2(new_n912), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n729), .A2(G330), .A3(new_n812), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n902), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT117), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n729), .A2(new_n902), .A3(new_n812), .A4(G330), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n815), .A2(new_n809), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1076), .A2(new_n1077), .A3(KEYINPUT117), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n811), .A2(new_n323), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n809), .B1(new_n703), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1078), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT118), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1078), .A2(new_n1086), .A3(KEYINPUT118), .A4(new_n1080), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1084), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1075), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n890), .A2(new_n894), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n903), .A2(new_n895), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(KEYINPUT116), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT116), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n903), .A2(new_n1096), .A3(new_n895), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n888), .B(new_n895), .C1(new_n1086), .C2(new_n1077), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1098), .A2(new_n1080), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1080), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1092), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1092), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n683), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n741), .B1(new_n275), .B2(new_n820), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n778), .A2(new_n310), .B1(new_n766), .B2(new_n215), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G116), .B2(new_n780), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n759), .A2(new_n770), .B1(new_n758), .B2(new_n202), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n251), .B(new_n1109), .C1(G87), .C2(new_n763), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n789), .A2(G294), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n1058), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n780), .A2(G132), .B1(new_n795), .B2(G128), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT119), .Z(new_n1114));
  NAND2_X1  g0914(.A1(new_n763), .A2(G150), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1115), .A2(KEYINPUT53), .B1(new_n797), .B2(new_n773), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(KEYINPUT53), .B2(new_n1115), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n789), .A2(G125), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n758), .A2(new_n208), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n251), .B1(new_n766), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G137), .C2(new_n777), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1112), .B1(new_n1114), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n746), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1106), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1093), .B2(new_n743), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n734), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1105), .A2(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1131), .A2(new_n781), .B1(new_n778), .B2(new_n836), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G125), .A2(new_n795), .B1(new_n767), .B2(G137), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n762), .B2(new_n1120), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G150), .C2(new_n774), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT59), .Z(new_n1136));
  AOI211_X1 g0936(.A(G33), .B(G41), .C1(new_n792), .C2(G159), .ZN(new_n1137));
  INV_X1    g0937(.A(G124), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n788), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT120), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n248), .A2(new_n259), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n577), .B2(new_n767), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n210), .B2(new_n770), .C1(new_n788), .C2(new_n759), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n215), .A2(new_n778), .B1(new_n781), .B2(new_n310), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n201), .A2(new_n758), .B1(new_n762), .B2(new_n253), .ZN(new_n1146));
  NOR4_X1   g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n952), .A4(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1142), .B(new_n208), .C1(G33), .C2(G41), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n746), .B1(new_n1141), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n820), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n735), .C1(G50), .C2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n292), .A2(new_n852), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT55), .Z(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n620), .B2(new_n295), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n295), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n1158), .C1(new_n618), .C2(new_n619), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1156), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n619), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT87), .B1(new_n303), .B2(new_n306), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n295), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1158), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n620), .A2(new_n295), .A3(new_n1159), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1155), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1154), .B1(new_n1171), .B2(new_n743), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n897), .A2(new_n908), .A3(new_n909), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1170), .B1(new_n923), .B2(G330), .ZN(new_n1174));
  OAI211_X1 g0974(.A(G330), .B(new_n1170), .C1(new_n926), .C2(new_n928), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(G330), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1171), .B1(new_n929), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n910), .A3(new_n1175), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1172), .B1(new_n1181), .B2(new_n734), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1075), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1184), .B(new_n1185), .C1(new_n1102), .C2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1187), .A2(new_n683), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1092), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1186), .B1(new_n1128), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1174), .A2(new_n1176), .A3(new_n1173), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n910), .B1(new_n1179), .B2(new_n1175), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT122), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT123), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1194), .A2(KEYINPUT123), .A3(new_n683), .A4(new_n1187), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1181), .B1(new_n1102), .B2(new_n1186), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1183), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1182), .B1(new_n1195), .B2(new_n1199), .ZN(G375));
  NOR2_X1   g1000(.A1(new_n902), .A2(new_n744), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT124), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n742), .B1(G68), .B2(new_n1153), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n777), .A2(G116), .B1(new_n795), .B2(G294), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n215), .B2(new_n762), .C1(new_n940), .C2(new_n788), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n780), .A2(G283), .B1(G107), .B2(new_n767), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1024), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1206), .A2(new_n248), .A3(new_n950), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1120), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n777), .A2(new_n1209), .B1(new_n795), .B2(G132), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n797), .B2(new_n762), .C1(new_n1131), .C2(new_n788), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n780), .A2(G137), .B1(G150), .B2(new_n767), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n248), .B1(new_n792), .B2(G58), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n208), .C2(new_n773), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1205), .A2(new_n1208), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1203), .B1(new_n746), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1091), .A2(new_n734), .B1(new_n1202), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1189), .A2(new_n985), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1075), .A2(new_n1091), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(G381));
  NAND3_X1  g1022(.A1(new_n1013), .A2(new_n807), .A3(new_n1044), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(G390), .A2(G384), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1009), .A2(new_n1224), .A3(new_n1221), .ZN(new_n1225));
  OR3_X1    g1025(.A1(new_n1225), .A2(G375), .A3(G378), .ZN(G407));
  INV_X1    g1026(.A(G378), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n659), .A2(G213), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G407), .B(G213), .C1(G375), .C2(new_n1230), .ZN(G409));
  NAND2_X1  g1031(.A1(G393), .A2(G396), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G390), .B1(new_n1232), .B2(new_n1223), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G390), .A2(new_n1232), .A3(new_n1223), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1234), .A2(new_n1009), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1009), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G378), .B(new_n1182), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1182), .B1(new_n1197), .B2(new_n985), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1227), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT125), .B1(new_n1075), .B2(new_n1091), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1244), .B(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n683), .A3(new_n1092), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1217), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n842), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(G384), .A3(new_n1217), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1242), .A2(new_n1243), .A3(new_n1228), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1229), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1228), .A2(KEYINPUT126), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1249), .A2(new_n1250), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1229), .A2(G2897), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1257), .B(new_n1258), .Z(new_n1259));
  OAI211_X1 g1059(.A(new_n1253), .B(new_n1254), .C1(new_n1255), .C2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1255), .B2(new_n1252), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1238), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1255), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1251), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1257), .B(new_n1258), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1264), .A2(new_n1267), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(G405));
  NAND2_X1  g1072(.A1(G375), .A2(new_n1227), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1239), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(new_n1252), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1252), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1238), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1275), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1264), .A2(new_n1279), .A3(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(G402));
endmodule


