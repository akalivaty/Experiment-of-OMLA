//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  AND2_X1   g000(.A1(KEYINPUT64), .A2(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT64), .A2(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(G146), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n187), .A2(new_n188), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(new_n195), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n194), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT66), .A3(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n209), .A3(new_n207), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT64), .A2(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n195), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n196), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n200), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n194), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n203), .A2(new_n214), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT30), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n210), .A2(G131), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(G128), .B1(new_n191), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n189), .A2(new_n226), .A3(G128), .A4(new_n192), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n205), .B2(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n208), .A2(KEYINPUT67), .A3(G134), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n207), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n223), .A2(new_n224), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n210), .B(new_n212), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n238), .B2(new_n202), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n214), .A2(new_n220), .A3(new_n240), .A4(new_n194), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n239), .A2(new_n241), .B1(new_n235), .B2(new_n230), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n237), .B1(new_n242), .B2(new_n224), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(G116), .B(G119), .Z(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT68), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT68), .B1(new_n247), .B2(new_n249), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT70), .B1(new_n243), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT72), .B(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(G210), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n258), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n238), .A2(new_n202), .A3(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n215), .A2(new_n216), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n191), .B1(new_n265), .B2(G146), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n266), .A2(new_n193), .B1(new_n219), .B2(new_n200), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n240), .B1(new_n267), .B2(new_n214), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n252), .B(new_n236), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n252), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n256), .A2(new_n263), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n223), .A2(new_n236), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n253), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n236), .B(new_n252), .C1(new_n202), .C2(new_n238), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n262), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n274), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n242), .A2(new_n252), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n271), .B2(new_n272), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n280), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n269), .A2(new_n270), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT71), .B1(new_n242), .B2(new_n252), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n277), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n281), .B1(new_n293), .B2(KEYINPUT28), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT73), .B1(new_n294), .B2(new_n262), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n256), .A2(new_n296), .A3(new_n262), .A4(new_n273), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n239), .A2(new_n241), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n224), .B1(new_n298), .B2(new_n236), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n223), .A2(new_n224), .A3(new_n236), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n253), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n253), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n262), .A3(new_n273), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT31), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(new_n263), .C1(new_n278), .C2(new_n281), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n295), .A2(new_n297), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT32), .ZN(new_n310));
  NOR2_X1   g124(.A1(G472), .A2(G902), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n290), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(KEYINPUT74), .B(new_n290), .C1(new_n312), .C2(new_n313), .ZN(new_n317));
  INV_X1    g131(.A(G128), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n229), .B1(new_n319), .B2(new_n266), .ZN(new_n320));
  INV_X1    g134(.A(G104), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(new_n321), .B2(G107), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  INV_X1    g137(.A(G107), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G104), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(G107), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n322), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n324), .A2(G104), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n321), .A2(G107), .ZN(new_n330));
  OAI21_X1  g144(.A(G101), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT80), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n333), .B(G101), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n320), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n228), .A2(new_n332), .A3(new_n229), .A4(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n214), .ZN(new_n339));
  NOR2_X1   g153(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n338), .B(new_n214), .C1(KEYINPUT81), .C2(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT10), .B1(new_n320), .B2(new_n335), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n322), .A2(new_n325), .A3(new_n327), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n347), .A2(G101), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n267), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n228), .A2(new_n229), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n335), .A3(KEYINPUT10), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n346), .A2(new_n352), .A3(new_n238), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G110), .B(G140), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT79), .ZN(new_n358));
  INV_X1    g172(.A(G227), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n352), .A2(new_n354), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n214), .B1(new_n364), .B2(new_n345), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n355), .A3(new_n361), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G469), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n355), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n362), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n356), .B2(new_n362), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n284), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n284), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT9), .B(G234), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G221), .B1(new_n378), .B2(G902), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G475), .A2(G902), .ZN(new_n381));
  AND2_X1   g195(.A1(KEYINPUT72), .A2(G237), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT72), .A2(G237), .ZN(new_n383));
  OAI211_X1 g197(.A(G214), .B(new_n260), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n197), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n259), .A2(new_n190), .A3(G214), .A4(new_n260), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT18), .A4(G131), .ZN(new_n387));
  NOR2_X1   g201(.A1(G125), .A2(G140), .ZN(new_n388));
  AND2_X1   g202(.A1(KEYINPUT76), .A2(G125), .ZN(new_n389));
  NOR2_X1   g203(.A1(KEYINPUT76), .A2(G125), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n391), .B2(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G146), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n195), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT83), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n385), .B2(new_n386), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT84), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n401), .B(new_n398), .C1(new_n385), .C2(new_n386), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n387), .B(new_n396), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n386), .ZN(new_n404));
  INV_X1    g218(.A(G131), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n385), .A2(new_n386), .A3(G131), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT16), .ZN(new_n409));
  INV_X1    g223(.A(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n391), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(G146), .B(new_n411), .C1(new_n392), .C2(new_n409), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n394), .A2(KEYINPUT19), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n392), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n195), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n403), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G113), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n321), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g236(.A1(KEYINPUT76), .A2(G125), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT76), .A2(G125), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(G140), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n388), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n409), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT76), .B(G125), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n428), .A2(KEYINPUT16), .A3(G140), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n195), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n412), .A3(KEYINPUT77), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(new_n195), .C1(new_n427), .C2(new_n429), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n406), .A2(new_n435), .A3(new_n407), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n407), .A2(new_n435), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n420), .B(new_n403), .C1(new_n434), .C2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n422), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n422), .B2(new_n439), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT20), .B(new_n381), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n422), .A2(new_n439), .ZN(new_n445));
  INV_X1    g259(.A(new_n381), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n439), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n431), .A2(new_n433), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n437), .A3(new_n436), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n420), .B1(new_n450), .B2(new_n403), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n284), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G475), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n443), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n443), .A2(KEYINPUT86), .A3(new_n447), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n459));
  INV_X1    g273(.A(G119), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G116), .ZN(new_n461));
  OAI211_X1 g275(.A(G113), .B(new_n461), .C1(new_n248), .C2(new_n459), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n335), .A2(new_n247), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n350), .A2(new_n351), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n252), .ZN(new_n465));
  XOR2_X1   g279(.A(G110), .B(G122), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n466), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n468), .B(new_n463), .C1(new_n464), .C2(new_n252), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n202), .A2(new_n391), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n228), .A2(new_n229), .A3(new_n428), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n473), .A2(G224), .A3(new_n260), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(G224), .B2(new_n260), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n465), .A2(new_n477), .A3(new_n466), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n474), .B1(new_n475), .B2(KEYINPUT7), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n462), .A2(new_n247), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n335), .B(new_n483), .Z(new_n484));
  XOR2_X1   g298(.A(new_n466), .B(KEYINPUT8), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n480), .A2(new_n469), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(new_n487), .A3(new_n284), .ZN(new_n488));
  OAI21_X1  g302(.A(G210), .B1(G237), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n479), .A2(new_n487), .A3(new_n284), .A4(new_n489), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n260), .A2(G952), .ZN(new_n494));
  NAND2_X1  g308(.A1(G234), .A2(G237), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT21), .B(G898), .Z(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(G902), .A3(G953), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT82), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G116), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(G122), .ZN(new_n505));
  INV_X1    g319(.A(G122), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT87), .B1(new_n506), .B2(G116), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n504), .A3(G122), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n324), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n511), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(G107), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n318), .A2(G143), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT89), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n205), .A2(KEYINPUT13), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n318), .B2(new_n197), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(G134), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  OAI21_X1  g338(.A(G107), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n510), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n522), .B(new_n205), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n513), .A2(new_n516), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G217), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n378), .A2(new_n532), .A3(G953), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n527), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n284), .ZN(new_n538));
  INV_X1    g352(.A(G478), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n540), .ZN(new_n541));
  NOR4_X1   g355(.A1(new_n380), .A2(new_n458), .A3(new_n503), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n532), .B1(G234), .B2(new_n284), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n318), .A2(G119), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n546), .A2(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n460), .A2(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(KEYINPUT23), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n548), .A2(new_n545), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT24), .B(G110), .Z(new_n552));
  OAI22_X1  g366(.A1(new_n550), .A2(G110), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n412), .A3(new_n395), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(G110), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n431), .A2(new_n555), .A3(new_n556), .A4(new_n433), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT22), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G137), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n554), .B(new_n564), .C1(new_n559), .C2(new_n560), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n284), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT25), .A4(new_n284), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n544), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n568), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n572), .B1(new_n544), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n316), .A2(new_n317), .A3(new_n542), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT90), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(new_n326), .ZN(G3));
  INV_X1    g391(.A(new_n536), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n535), .B1(new_n527), .B2(new_n530), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT33), .B1(new_n534), .B2(new_n536), .ZN(new_n582));
  OAI21_X1  g396(.A(G478), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n537), .A2(new_n539), .A3(new_n284), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n539), .A2(new_n284), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n456), .B2(new_n457), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n503), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT91), .Z(new_n591));
  NAND2_X1  g405(.A1(new_n309), .A2(new_n284), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n309), .A2(new_n311), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n380), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n574), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NOR2_X1   g415(.A1(new_n441), .A2(new_n442), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n444), .B1(new_n602), .B2(new_n446), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n603), .A2(new_n453), .A3(new_n443), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n541), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n597), .A2(new_n503), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT35), .B(G107), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT92), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n606), .B(new_n608), .ZN(G9));
  NAND2_X1  g423(.A1(new_n570), .A2(new_n571), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n543), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n565), .A2(KEYINPUT36), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n561), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n561), .A2(new_n613), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n543), .A2(G902), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT93), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n458), .A2(new_n503), .A3(new_n541), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n596), .A2(new_n620), .A3(new_n595), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT37), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G110), .ZN(G12));
  NAND4_X1  g438(.A1(new_n316), .A2(new_n620), .A3(new_n317), .A4(new_n596), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n496), .B1(new_n498), .B2(G900), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n604), .A2(new_n541), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n493), .A2(new_n502), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(KEYINPUT94), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n627), .B2(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n625), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n318), .ZN(G30));
  XNOR2_X1  g451(.A(new_n626), .B(KEYINPUT39), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n596), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT40), .Z(new_n640));
  NOR2_X1   g454(.A1(new_n572), .A2(new_n617), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n263), .B1(new_n256), .B2(new_n273), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n286), .B2(new_n263), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n312), .B2(new_n313), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n458), .ZN(new_n648));
  INV_X1    g462(.A(new_n541), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n493), .B(KEYINPUT38), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n647), .A2(new_n502), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n197), .ZN(G45));
  NAND2_X1  g467(.A1(new_n594), .A2(KEYINPUT32), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT74), .B1(new_n656), .B2(new_n290), .ZN(new_n657));
  INV_X1    g471(.A(new_n317), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT95), .ZN(new_n660));
  INV_X1    g474(.A(new_n587), .ZN(new_n661));
  AND4_X1   g475(.A1(new_n660), .A2(new_n458), .A3(new_n661), .A4(new_n626), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n660), .B1(new_n588), .B2(new_n626), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n662), .A2(new_n663), .A3(new_n629), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n659), .A2(new_n596), .A3(new_n620), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  NAND2_X1  g480(.A1(new_n371), .A2(new_n284), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n373), .ZN(new_n669));
  INV_X1    g483(.A(new_n379), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n316), .A2(new_n317), .A3(new_n574), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n591), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT41), .B(G113), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NOR2_X1   g489(.A1(new_n605), .A2(new_n503), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  AND4_X1   g492(.A1(new_n316), .A2(new_n620), .A3(new_n317), .A4(new_n671), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n621), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  NAND2_X1  g495(.A1(new_n287), .A2(new_n263), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n297), .A2(new_n306), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n311), .B(KEYINPUT96), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT97), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n592), .B2(G472), .ZN(new_n687));
  INV_X1    g501(.A(G472), .ZN(new_n688));
  AOI211_X1 g502(.A(KEYINPUT97), .B(new_n688), .C1(new_n309), .C2(new_n284), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n574), .B(new_n685), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n650), .A2(new_n671), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n690), .A2(new_n503), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n506), .ZN(G24));
  OAI211_X1 g507(.A(new_n619), .B(new_n685), .C1(new_n687), .C2(new_n689), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n458), .A2(new_n661), .A3(new_n626), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT95), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n588), .A2(new_n660), .A3(new_n626), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(KEYINPUT98), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n662), .B2(new_n663), .ZN(new_n701));
  INV_X1    g515(.A(new_n671), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n629), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n695), .A2(new_n699), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n363), .A2(KEYINPUT99), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT99), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n356), .A2(new_n708), .A3(new_n362), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(G469), .A3(new_n709), .A4(new_n366), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT100), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n708), .B1(new_n356), .B2(new_n362), .ZN(new_n712));
  AOI211_X1 g526(.A(KEYINPUT99), .B(new_n361), .C1(new_n344), .C2(new_n355), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n715), .A3(G469), .A4(new_n366), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n711), .A2(new_n716), .A3(new_n373), .A4(new_n375), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n379), .ZN(new_n718));
  INV_X1    g532(.A(new_n493), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n502), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n316), .A2(new_n317), .A3(new_n574), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n701), .A2(new_n699), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n706), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n314), .A2(new_n574), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n706), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n699), .A3(new_n701), .A4(new_n721), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT101), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  AND4_X1   g544(.A1(new_n316), .A2(new_n317), .A3(new_n574), .A4(new_n721), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n628), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  OR2_X1    g547(.A1(new_n367), .A2(KEYINPUT45), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n366), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(G469), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT46), .B1(new_n736), .B2(new_n375), .ZN(new_n737));
  INV_X1    g551(.A(new_n373), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n375), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n670), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n638), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT102), .Z(new_n743));
  NAND2_X1  g557(.A1(new_n648), .A2(new_n661), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n595), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n619), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n720), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n743), .B(new_n750), .C1(new_n749), .C2(new_n748), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  XNOR2_X1  g566(.A(new_n741), .B(KEYINPUT47), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n574), .A2(new_n720), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n621), .A2(new_n679), .B1(new_n672), .B2(new_n676), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n692), .B1(new_n591), .B2(new_n672), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n759), .A2(new_n728), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n316), .A2(new_n620), .A3(new_n317), .A4(new_n596), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n720), .A2(new_n541), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n604), .A3(new_n626), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n648), .A2(new_n541), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n597), .A2(new_n503), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n622), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n595), .A2(new_n590), .A3(new_n574), .A4(new_n596), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n575), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n575), .B2(new_n771), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n766), .B(new_n769), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n701), .A2(new_n699), .A3(new_n721), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n695), .A2(new_n777), .B1(new_n731), .B2(new_n628), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n759), .A2(new_n728), .A3(new_n760), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n763), .A2(new_n776), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n764), .A2(new_n634), .ZN(new_n782));
  INV_X1    g596(.A(new_n626), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT105), .B1(new_n619), .B2(new_n783), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n572), .A2(new_n617), .A3(KEYINPUT105), .A4(new_n783), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n718), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT106), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n648), .A2(new_n629), .A3(new_n649), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n646), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n646), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n373), .A2(new_n375), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(KEYINPUT100), .B2(new_n710), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n670), .B1(new_n793), .B2(new_n716), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT105), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n641), .B2(new_n626), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n796), .B2(new_n785), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT106), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n782), .A2(new_n665), .A3(new_n704), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT107), .B1(new_n800), .B2(new_n801), .ZN(new_n805));
  INV_X1    g619(.A(new_n664), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n592), .A2(new_n686), .A3(G472), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n619), .A3(new_n685), .A4(new_n703), .ZN(new_n810));
  OAI22_X1  g624(.A1(new_n625), .A2(new_n806), .B1(new_n723), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n636), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT52), .A4(new_n799), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n800), .A2(KEYINPUT108), .A3(new_n801), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n804), .A2(new_n805), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n805), .A2(new_n814), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n800), .A2(KEYINPUT108), .A3(new_n801), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT108), .B1(new_n800), .B2(new_n801), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n781), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT104), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n776), .A2(new_n761), .A3(new_n825), .A4(new_n778), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n575), .A2(new_n771), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT103), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n772), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n769), .A3(new_n766), .A4(new_n778), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT104), .B1(new_n830), .B2(new_n779), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n800), .B(new_n801), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(new_n758), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n824), .A2(new_n834), .A3(KEYINPUT54), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n826), .A2(new_n831), .A3(KEYINPUT53), .A4(new_n832), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT111), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n822), .B1(new_n818), .B2(new_n821), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n826), .A2(new_n831), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT110), .B(new_n758), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n817), .B2(new_n823), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(KEYINPUT53), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n838), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n836), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n656), .A2(new_n574), .A3(new_n645), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n702), .A2(new_n496), .A3(new_n720), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n588), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n746), .A2(new_n852), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT115), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n695), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n851), .A2(new_n648), .A3(new_n587), .A4(new_n852), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n746), .A2(new_n495), .A3(new_n494), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n690), .ZN(new_n860));
  INV_X1    g674(.A(new_n651), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n501), .A3(new_n861), .A4(new_n671), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(KEYINPUT114), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n862), .B2(KEYINPUT114), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n857), .B(new_n858), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n669), .A2(new_n379), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n753), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n720), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n854), .B(KEYINPUT51), .C1(new_n867), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n866), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n864), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n871), .A3(new_n857), .A4(new_n858), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT51), .B1(new_n877), .B2(new_n854), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n494), .B(new_n853), .C1(new_n874), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n725), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n856), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT48), .Z(new_n882));
  NOR4_X1   g696(.A1(new_n859), .A2(new_n629), .A3(new_n702), .A4(new_n690), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n849), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n669), .B(KEYINPUT49), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n886), .A2(new_n651), .A3(new_n670), .A4(new_n501), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n851), .A2(new_n887), .A3(new_n648), .A4(new_n661), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(G75));
  INV_X1    g703(.A(new_n781), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n839), .B2(new_n840), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n833), .A2(new_n758), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n284), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G210), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n470), .A2(new_n478), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n476), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(KEYINPUT56), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n894), .B2(new_n895), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n260), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n375), .A2(KEYINPUT57), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n848), .B1(new_n891), .B2(new_n892), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n835), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n375), .A2(KEYINPUT57), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n371), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n736), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n893), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n904), .B1(new_n910), .B2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(new_n602), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n602), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n904), .ZN(G60));
  INV_X1    g731(.A(new_n904), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n585), .B(KEYINPUT59), .Z(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n907), .B2(new_n835), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n581), .A2(new_n582), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n849), .A2(new_n919), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n922), .ZN(G63));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT118), .Z(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n891), .B2(new_n892), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n614), .A2(new_n615), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n566), .A2(new_n567), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n935), .B2(new_n931), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n926), .B1(new_n936), .B2(new_n904), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n824), .B2(new_n834), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n939), .A2(KEYINPUT119), .A3(new_n934), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT119), .B1(new_n939), .B2(new_n934), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n918), .A2(KEYINPUT61), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n931), .B2(new_n932), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n931), .B2(new_n935), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n939), .A2(KEYINPUT119), .A3(new_n934), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n938), .A2(new_n947), .A3(new_n944), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n937), .B1(new_n945), .B2(new_n949), .ZN(G66));
  AOI21_X1  g764(.A(new_n260), .B1(new_n497), .B2(G224), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n829), .A2(new_n769), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n759), .A2(new_n760), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n955), .B2(new_n260), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT121), .B(KEYINPUT122), .Z(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(G898), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n896), .B1(new_n959), .B2(G953), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  XOR2_X1   g775(.A(new_n415), .B(KEYINPUT123), .Z(new_n962));
  XNOR2_X1  g776(.A(new_n243), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(G900), .A2(G953), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n751), .A2(new_n756), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n812), .A2(new_n728), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n743), .A2(new_n880), .A3(new_n789), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(new_n732), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n963), .B(new_n964), .C1(new_n968), .C2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n652), .A2(new_n812), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n767), .A2(new_n589), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n639), .A2(new_n720), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n659), .A2(new_n574), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n965), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n969), .B1(new_n979), .B2(new_n963), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT126), .B1(new_n979), .B2(new_n963), .ZN(new_n981));
  INV_X1    g795(.A(G900), .ZN(new_n982));
  OAI21_X1  g796(.A(G953), .B1(new_n359), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT125), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n980), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  OAI221_X1 g800(.A(new_n969), .B1(KEYINPUT126), .B2(new_n984), .C1(new_n979), .C2(new_n963), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G72));
  XNOR2_X1  g802(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n688), .A2(new_n284), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n968), .B2(new_n955), .ZN(new_n992));
  INV_X1    g806(.A(new_n274), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n991), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n978), .B2(new_n954), .ZN(new_n996));
  INV_X1    g810(.A(new_n642), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n994), .B(new_n918), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n847), .A2(new_n993), .A3(new_n995), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(G57));
endmodule


