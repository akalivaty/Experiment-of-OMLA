//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G68), .A2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G58), .C2(G232), .ZN(new_n220));
  INV_X1    g0020(.A(new_n206), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n210), .B(new_n223), .C1(new_n226), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n213), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n212), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n247));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(new_n247), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G238), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n259), .A2(new_n260), .B1(new_n231), .B2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G226), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n256), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n250), .B(new_n254), .C1(new_n265), .C2(new_n252), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n264), .B1(G232), .B2(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n255), .ZN(new_n271));
  INV_X1    g0071(.A(new_n252), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(new_n250), .A4(new_n254), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT74), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n267), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n271), .A2(new_n272), .B1(G238), .B2(new_n253), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(KEYINPUT74), .A3(new_n274), .A4(new_n250), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G169), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT14), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n277), .A2(KEYINPUT14), .A3(G169), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n267), .ZN(new_n285));
  INV_X1    g0085(.A(new_n275), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n224), .B1(new_n206), .B2(new_n258), .ZN(new_n292));
  OR3_X1    g0092(.A1(new_n258), .A2(KEYINPUT68), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n225), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n225), .B2(G68), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G50), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n292), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT71), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n246), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(new_n292), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n246), .A2(G20), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT12), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G68), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n304), .A2(new_n308), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n284), .A2(new_n321), .A3(new_n289), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n291), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n285), .A2(new_n286), .A3(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n277), .A2(G200), .A3(new_n279), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n253), .A2(G244), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT3), .B(G33), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(G232), .A3(new_n263), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(G238), .A3(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G107), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n331), .B(new_n332), .C1(new_n333), .C2(new_n330), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n249), .B(new_n329), .C1(new_n334), .C2(new_n272), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT70), .B(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g0137(.A(KEYINPUT15), .B(G87), .Z(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n294), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n341), .A2(new_n300), .B1(new_n225), .B2(new_n297), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n292), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n312), .A2(new_n297), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n316), .C2(new_n297), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n337), .B(new_n345), .C1(G169), .C2(new_n335), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n323), .A2(new_n328), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT17), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n330), .B2(G20), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n268), .A2(new_n269), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n202), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G58), .A2(G68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(G58), .A3(G68), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n358), .A3(new_n203), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G20), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n299), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n349), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n352), .B2(new_n225), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n268), .A2(new_n269), .A3(new_n350), .A4(G20), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n359), .A2(G20), .B1(G159), .B2(new_n299), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(new_n368), .A3(new_n292), .ZN(new_n369));
  INV_X1    g0169(.A(new_n341), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n315), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n306), .A2(new_n292), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n371), .A2(new_n372), .B1(new_n306), .B2(new_n341), .ZN(new_n373));
  OAI211_X1 g0173(.A(G226), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n330), .A2(KEYINPUT77), .A3(G226), .A4(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n330), .A2(G223), .A3(new_n263), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT78), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n272), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT81), .B(G190), .Z(new_n385));
  INV_X1    g0185(.A(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n252), .A2(new_n247), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n231), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n252), .A2(new_n247), .A3(KEYINPUT79), .A4(G232), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n249), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(G200), .B1(new_n384), .B2(new_n390), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n369), .B(new_n373), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT82), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n348), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n392), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n369), .A2(new_n373), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT82), .A4(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n369), .A2(new_n373), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n384), .A2(new_n336), .A3(new_n390), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(G169), .B1(new_n384), .B2(new_n390), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT80), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n384), .A2(new_n390), .ZN(new_n408));
  INV_X1    g0208(.A(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT80), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n406), .B1(new_n404), .B2(new_n405), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .A3(new_n402), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n401), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(KEYINPUT66), .A2(G223), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT66), .A2(G223), .ZN(new_n421));
  OAI21_X1  g0221(.A(G1698), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n263), .A2(G222), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n330), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n272), .C1(G77), .C2(new_n330), .ZN(new_n425));
  OR2_X1    g0225(.A1(KEYINPUT65), .A2(G226), .ZN(new_n426));
  NAND2_X1  g0226(.A1(KEYINPUT65), .A2(G226), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n253), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n250), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT67), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT67), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n425), .A2(new_n431), .A3(new_n250), .A4(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G190), .ZN(new_n434));
  INV_X1    g0234(.A(G150), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n296), .A2(new_n341), .B1(new_n435), .B2(new_n300), .ZN(new_n436));
  INV_X1    g0236(.A(new_n203), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n225), .B1(new_n437), .B2(new_n301), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n292), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT9), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n306), .A2(new_n301), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n315), .A2(G50), .A3(new_n372), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n439), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n341), .B1(new_n293), .B2(new_n295), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n300), .A2(new_n435), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n444), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n292), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n441), .B(new_n442), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT9), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n430), .A2(G200), .A3(new_n432), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n434), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n433), .A2(G190), .B1(KEYINPUT73), .B2(KEYINPUT10), .ZN(new_n456));
  INV_X1    g0256(.A(new_n454), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n450), .A4(new_n451), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n448), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n433), .B2(new_n336), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(G169), .B2(new_n433), .ZN(new_n463));
  INV_X1    g0263(.A(G200), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n335), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT72), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n345), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n335), .A2(G190), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n345), .A2(new_n466), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n419), .A2(new_n460), .A3(new_n463), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n347), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n212), .B1(new_n246), .B2(G33), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n313), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT86), .B(G116), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n312), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n225), .C1(G33), .C2(new_n217), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n292), .B(new_n479), .C1(new_n475), .C2(new_n225), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT20), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n474), .B(new_n477), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G264), .A2(G1698), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n330), .B(new_n485), .C1(new_n218), .C2(G1698), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n272), .C1(G303), .C2(new_n330), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  INV_X1    g0290(.A(new_n224), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n488), .A2(new_n490), .B1(new_n491), .B2(new_n251), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G270), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(G274), .A3(new_n490), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n487), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n484), .A2(new_n495), .A3(G169), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n495), .A2(new_n287), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n484), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n484), .A2(new_n495), .A3(KEYINPUT21), .A4(G169), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n484), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n495), .A2(new_n385), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(G200), .B2(new_n495), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT22), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n212), .A2(KEYINPUT86), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT86), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n510), .A3(G33), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n225), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n330), .A2(new_n225), .A3(G87), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n225), .A2(G107), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT23), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n512), .A2(new_n225), .B1(new_n514), .B2(new_n515), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n518), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n292), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n372), .B1(G1), .B2(new_n258), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n333), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n306), .A2(new_n333), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n529), .B(KEYINPUT25), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n525), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n533));
  OAI211_X1 g0333(.A(G250), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G294), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n272), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n492), .A2(G264), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n494), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G190), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n537), .A2(KEYINPUT88), .A3(new_n538), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT88), .B1(new_n537), .B2(new_n538), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n494), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(new_n464), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n532), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n447), .B1(new_n520), .B2(new_n523), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n527), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(G169), .ZN(new_n548));
  OAI211_X1 g0348(.A(G179), .B(new_n494), .C1(new_n541), .C2(new_n542), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(new_n531), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT83), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT6), .ZN(new_n553));
  AND2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n333), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n225), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n300), .A2(new_n297), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n552), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n559), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n333), .A2(KEYINPUT6), .A3(G97), .ZN(new_n562));
  XNOR2_X1  g0362(.A(G97), .B(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n553), .ZN(new_n564));
  OAI211_X1 g0364(.A(KEYINPUT83), .B(new_n561), .C1(new_n564), .C2(new_n225), .ZN(new_n565));
  OAI21_X1  g0365(.A(G107), .B1(new_n364), .B2(new_n365), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n292), .B1(new_n217), .B2(new_n306), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT84), .B1(new_n492), .B2(G257), .ZN(new_n569));
  AND2_X1   g0369(.A1(KEYINPUT5), .A2(G41), .ZN(new_n570));
  NOR2_X1   g0370(.A1(KEYINPUT5), .A2(G41), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n490), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND4_X1   g0372(.A1(KEYINPUT84), .A2(new_n572), .A3(G257), .A4(new_n252), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n494), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n330), .A2(G244), .A3(new_n263), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(G33), .B2(G283), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .ZN(new_n578));
  INV_X1    g0378(.A(G250), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n263), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n330), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n252), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(G200), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n575), .A2(new_n576), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n478), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n272), .ZN(new_n586));
  INV_X1    g0386(.A(new_n494), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n492), .A2(KEYINPUT84), .A3(G257), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n572), .A2(G257), .A3(new_n252), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n587), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n592), .A3(G190), .ZN(new_n593));
  INV_X1    g0393(.A(new_n526), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G97), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n568), .A2(new_n583), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n338), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n225), .B1(new_n255), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n555), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n225), .A2(G33), .A3(G97), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n599), .A2(new_n601), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n330), .A2(new_n225), .A3(G68), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n292), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n338), .B1(new_n310), .B2(new_n311), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT87), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n447), .B1(new_n603), .B2(new_n604), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n610), .A2(new_n611), .A3(new_n607), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n597), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n252), .B(G250), .C1(G1), .C2(new_n489), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n330), .A2(G244), .A3(G1698), .ZN(new_n616));
  OAI211_X1 g0416(.A(G238), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n511), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n615), .B1(new_n618), .B2(new_n272), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n490), .A2(G274), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n409), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n336), .A3(new_n620), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n613), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n606), .A2(KEYINPUT87), .A3(new_n608), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n611), .B1(new_n610), .B2(new_n607), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n625), .A2(new_n626), .B1(G87), .B2(new_n594), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n464), .B1(new_n619), .B2(new_n620), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n619), .A2(G190), .A3(new_n620), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n596), .A2(new_n624), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n567), .A2(new_n292), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n306), .A2(new_n217), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(new_n595), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n568), .B2(new_n595), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(G169), .B1(new_n586), .B2(new_n592), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n574), .A2(new_n582), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n336), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n632), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n472), .A2(new_n506), .A3(new_n551), .A4(new_n643), .ZN(G372));
  INV_X1    g0444(.A(new_n463), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n402), .A2(new_n403), .A3(new_n410), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(new_n413), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n327), .A2(new_n346), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n321), .B1(new_n284), .B2(new_n289), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT75), .B(new_n288), .C1(new_n282), .C2(new_n283), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n651), .B2(new_n320), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n647), .B1(new_n652), .B2(new_n401), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n645), .B1(new_n653), .B2(new_n460), .ZN(new_n654));
  INV_X1    g0454(.A(new_n472), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n624), .B(KEYINPUT89), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n635), .A2(KEYINPUT85), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n568), .A2(new_n637), .A3(new_n595), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n642), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n624), .A2(new_n631), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT26), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n537), .A2(new_n538), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n537), .A2(KEYINPUT88), .A3(new_n538), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(G200), .B1(new_n666), .B2(new_n494), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n547), .B(new_n531), .C1(new_n667), .C2(new_n540), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n550), .B2(new_n502), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n625), .A2(new_n626), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(new_n597), .B1(new_n409), .B2(new_n621), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n619), .A2(G190), .A3(new_n620), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n628), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n671), .A2(new_n623), .B1(new_n673), .B2(new_n627), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n659), .A2(new_n674), .A3(new_n596), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n656), .B(new_n661), .C1(new_n669), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n641), .A2(new_n336), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(G169), .B2(new_n641), .ZN(new_n678));
  INV_X1    g0478(.A(new_n635), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n674), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n654), .B1(new_n655), .B2(new_n684), .ZN(G369));
  NAND2_X1  g0485(.A1(new_n549), .A2(new_n548), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n532), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n668), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G13), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G20), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n246), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n688), .B1(new_n532), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n550), .B2(new_n696), .ZN(new_n698));
  INV_X1    g0498(.A(new_n696), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n502), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n503), .A2(new_n699), .ZN(new_n702));
  MUX2_X1   g0502(.A(new_n506), .B(new_n502), .S(new_n702), .Z(new_n703));
  NOR2_X1   g0503(.A1(new_n688), .A2(new_n700), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n701), .A2(G330), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n502), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n545), .B1(new_n707), .B2(new_n687), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n699), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n207), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n601), .A2(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n227), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(new_n699), .C1(new_n676), .C2(new_n682), .ZN(new_n719));
  INV_X1    g0519(.A(new_n656), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n708), .B2(new_n643), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT26), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n680), .B2(new_n674), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n659), .A2(new_n660), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n696), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n726), .B2(new_n718), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n643), .A2(new_n551), .A3(new_n506), .A4(new_n699), .ZN(new_n729));
  INV_X1    g0529(.A(new_n621), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n666), .A2(new_n641), .A3(new_n499), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n495), .A2(new_n336), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n586), .A2(new_n592), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n543), .A2(new_n735), .A3(new_n736), .A4(new_n621), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n696), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n728), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n717), .B1(new_n745), .B2(G1), .ZN(G364));
  OR2_X1    g0546(.A1(new_n703), .A2(G330), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT90), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n703), .A2(G330), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n246), .B1(new_n690), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n712), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n748), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n224), .B1(G20), .B2(new_n409), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n336), .A2(new_n225), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n385), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n324), .A3(new_n464), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G326), .A2(new_n759), .B1(new_n761), .B2(G311), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n324), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n225), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT93), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n225), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(new_n324), .A3(new_n464), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(G329), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n324), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  INV_X1    g0573(.A(G303), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n352), .B1(new_n772), .B2(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n757), .A2(new_n464), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n385), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n771), .B(new_n776), .C1(G322), .C2(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n758), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI221_X1 g0583(.A(new_n780), .B1(KEYINPUT93), .B2(new_n766), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n759), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n301), .A2(new_n785), .B1(new_n782), .B2(new_n202), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n765), .A2(new_n217), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT32), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n769), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n333), .B2(new_n772), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n790), .A2(new_n788), .B1(new_n600), .B2(new_n775), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n786), .A2(new_n352), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n778), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n760), .A2(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n760), .A2(KEYINPUT92), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n794), .B1(new_n201), .B2(new_n795), .C1(new_n297), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n756), .B1(new_n784), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n755), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n241), .A2(G45), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n711), .A2(new_n330), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(G45), .C2(new_n227), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n330), .A2(new_n207), .ZN(new_n808));
  XNOR2_X1  g0608(.A(G355), .B(KEYINPUT91), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(G116), .B2(new_n207), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n800), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n803), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n752), .C1(new_n703), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n754), .A2(new_n813), .ZN(G396));
  NOR2_X1   g0614(.A1(new_n346), .A2(new_n696), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n345), .A2(new_n696), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n470), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n817), .B2(new_n346), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n699), .B(new_n818), .C1(new_n676), .C2(new_n682), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT96), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n743), .B(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n818), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n684), .B2(new_n696), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n822), .B(new_n824), .Z(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n753), .ZN(new_n826));
  INV_X1    g0626(.A(new_n772), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G68), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n301), .B2(new_n775), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT95), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(KEYINPUT95), .ZN(new_n831));
  INV_X1    g0631(.A(new_n765), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n352), .B1(new_n832), .B2(G58), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G137), .A2(new_n759), .B1(new_n781), .B2(G150), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT94), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n795), .C1(new_n789), .C2(new_n798), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  AOI211_X1 g0639(.A(new_n834), .B(new_n839), .C1(G132), .C2(new_n770), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n785), .A2(new_n774), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n772), .A2(new_n600), .ZN(new_n842));
  INV_X1    g0642(.A(new_n775), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n787), .C1(G107), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n778), .A2(G294), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n781), .A2(G283), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n330), .B1(new_n770), .B2(G311), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n798), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n841), .B(new_n848), .C1(new_n475), .C2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n755), .B1(new_n840), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n823), .A2(new_n801), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n755), .A2(new_n801), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n297), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n851), .A2(new_n752), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n826), .A2(new_n855), .ZN(G384));
  AOI21_X1  g0656(.A(KEYINPUT37), .B1(new_n398), .B2(new_n399), .ZN(new_n857));
  INV_X1    g0657(.A(new_n694), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n402), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n412), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n646), .A2(new_n393), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT98), .B1(new_n402), .B2(new_n858), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n863), .B(new_n694), .C1(new_n369), .C2(new_n373), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n862), .A2(new_n864), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n867), .B(KEYINPUT38), .C1(new_n419), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n395), .A2(new_n400), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n859), .B1(new_n871), .B2(new_n647), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n402), .B1(new_n417), .B2(new_n858), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n646), .A2(new_n393), .A3(new_n859), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(new_n857), .B1(KEYINPUT37), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n870), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT101), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n740), .A2(new_n741), .A3(new_n818), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n320), .A2(new_n696), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n323), .A2(new_n328), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n320), .B(new_n696), .C1(new_n651), .C2(new_n327), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n414), .A2(new_n418), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n868), .B1(new_n888), .B2(new_n871), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n868), .A2(new_n393), .A3(new_n646), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .B1(new_n857), .B2(new_n873), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n870), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n869), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n885), .A2(new_n884), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(new_n742), .A3(new_n894), .A4(new_n818), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n742), .A2(new_n472), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n898), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT99), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n323), .B2(new_n696), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n651), .A2(KEYINPUT99), .A3(new_n320), .A4(new_n699), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n892), .B2(new_n869), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n869), .A2(new_n876), .A3(new_n906), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT100), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n869), .A2(new_n876), .A3(new_n906), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT100), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n905), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n815), .B(KEYINPUT97), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n819), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n894), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n869), .B2(new_n892), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n647), .A2(new_n858), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n913), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n727), .A2(new_n472), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n654), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n901), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n246), .B2(new_n690), .ZN(new_n924));
  INV_X1    g0724(.A(new_n564), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n212), .B1(new_n925), .B2(KEYINPUT35), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n226), .C1(KEYINPUT35), .C2(new_n925), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n228), .A2(G77), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n356), .A2(new_n358), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n929), .A2(new_n930), .B1(G50), .B2(new_n202), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n689), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n924), .A2(new_n928), .A3(new_n932), .ZN(G367));
  NOR2_X1   g0733(.A1(new_n627), .A2(new_n699), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n660), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n720), .B2(new_n934), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT43), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n659), .B(new_n596), .C1(new_n679), .C2(new_n699), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT102), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n680), .A2(new_n696), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n659), .B1(new_n943), .B2(new_n687), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT103), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n699), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n704), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT42), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n938), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n936), .A2(new_n937), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n706), .A2(new_n943), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT104), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n952), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n955), .ZN(new_n958));
  INV_X1    g0758(.A(new_n956), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n951), .A2(new_n952), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n712), .B(KEYINPUT41), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n942), .A2(new_n709), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n709), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n940), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT109), .A3(new_n706), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n706), .A2(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n706), .A2(KEYINPUT109), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n967), .A2(new_n974), .A3(new_n975), .A4(new_n971), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n701), .A2(new_n705), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n749), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n979), .A2(new_n706), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n745), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT108), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT107), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n745), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n983), .B1(new_n982), .B2(new_n985), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n963), .B1(new_n989), .B2(new_n745), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n957), .B(new_n961), .C1(new_n990), .C2(new_n751), .ZN(new_n991));
  INV_X1    g0791(.A(new_n806), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n804), .B1(new_n207), .B2(new_n339), .C1(new_n237), .C2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(G317), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n352), .B1(new_n769), .B2(new_n994), .C1(new_n765), .C2(new_n333), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n843), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT46), .B1(new_n843), .B2(new_n475), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n772), .A2(new_n217), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G294), .A2(new_n781), .B1(new_n759), .B2(G311), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n798), .C2(new_n773), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G303), .B2(new_n778), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n352), .B1(new_n843), .B2(G58), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n832), .A2(G68), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n297), .C2(new_n772), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G143), .B2(new_n759), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n798), .A2(new_n301), .B1(new_n789), .B2(new_n782), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT110), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1006), .B1(new_n435), .B2(new_n795), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n770), .A2(G137), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1002), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n752), .B(new_n993), .C1(new_n1013), .C2(new_n756), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT111), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n936), .A2(new_n803), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n991), .A2(new_n1018), .ZN(G387));
  AOI22_X1  g0819(.A1(G311), .A2(new_n781), .B1(new_n759), .B2(G322), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n774), .B2(new_n798), .C1(new_n994), .C2(new_n795), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n773), .B2(new_n765), .C1(new_n763), .C2(new_n775), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n770), .A2(G326), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n330), .B1(new_n827), .B2(new_n475), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n339), .A2(new_n765), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n778), .B2(G50), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT113), .Z(new_n1033));
  NOR2_X1   g0833(.A1(new_n782), .A2(new_n341), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n760), .A2(new_n202), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n330), .B1(new_n769), .B2(new_n435), .C1(new_n297), .C2(new_n775), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1034), .A2(new_n998), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n759), .A2(G159), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT112), .Z(new_n1039));
  NAND3_X1  g0839(.A1(new_n1033), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n756), .B1(new_n1030), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G116), .B(new_n601), .C1(G68), .C2(G77), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n341), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT50), .B1(new_n341), .B2(G50), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n489), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n992), .B1(new_n234), .B2(G45), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n808), .A2(new_n714), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n711), .A2(new_n333), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n803), .B(new_n755), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1041), .A2(new_n753), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT115), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n698), .A2(new_n803), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1052), .A2(new_n1053), .B1(new_n751), .B2(new_n980), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n982), .A2(new_n985), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n712), .C1(new_n745), .C2(new_n980), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(G393));
  INV_X1    g0857(.A(new_n1055), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n989), .B(new_n712), .C1(new_n977), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n977), .A2(new_n751), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G311), .A2(new_n778), .B1(new_n759), .B2(G317), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  AOI22_X1  g0862(.A1(G283), .A2(new_n843), .B1(new_n770), .B2(G322), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT116), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n782), .A2(new_n774), .B1(new_n333), .B2(new_n772), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n352), .B1(new_n765), .B2(new_n476), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1063), .A2(KEYINPUT116), .B1(new_n763), .B2(new_n760), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1062), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G150), .A2(new_n759), .B1(new_n778), .B2(G159), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n832), .A2(G77), .B1(new_n843), .B2(G68), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n837), .B2(new_n769), .C1(new_n782), .C2(new_n301), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n849), .B2(new_n370), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n330), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n1075), .B2(new_n842), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT117), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n753), .B1(new_n1077), .B2(new_n755), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n804), .B1(new_n217), .B2(new_n207), .C1(new_n244), .C2(new_n992), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n812), .C2(new_n942), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1059), .A2(new_n1060), .A3(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(KEYINPUT119), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n916), .A2(new_n905), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n909), .A2(new_n1083), .A3(new_n912), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n903), .A2(KEYINPUT118), .A3(new_n904), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT118), .B1(new_n903), .B2(new_n904), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  MUX2_X1   g0887(.A(new_n681), .B(new_n724), .S(new_n722), .Z(new_n1088));
  OAI21_X1  g0888(.A(new_n656), .B1(new_n669), .B2(new_n675), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n699), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n817), .A2(new_n346), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1090), .A2(new_n1092), .B1(new_n346), .B2(new_n696), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n894), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1087), .A2(new_n881), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n742), .A2(new_n894), .A3(G330), .A4(new_n818), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1084), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1084), .B2(new_n1095), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n742), .A2(new_n472), .A3(G330), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n920), .A2(new_n654), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n815), .B1(new_n726), .B2(new_n1091), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n740), .A2(new_n741), .A3(G330), .A4(new_n818), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n884), .A3(new_n885), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1096), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n915), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1096), .B2(new_n1103), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1100), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1097), .A2(new_n1098), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1082), .B1(new_n1108), .B2(new_n713), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1096), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1084), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n920), .A2(new_n654), .A3(new_n1099), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n915), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1113), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(KEYINPUT119), .A3(new_n712), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1109), .A2(new_n1110), .A3(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1097), .A2(new_n1098), .A3(new_n750), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n828), .B1(new_n600), .B2(new_n775), .C1(new_n297), .C2(new_n765), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n352), .B1(new_n763), .B2(new_n769), .C1(new_n795), .C2(new_n212), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(G107), .C2(new_n781), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n217), .B2(new_n798), .C1(new_n773), .C2(new_n785), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n330), .B1(new_n772), .B2(new_n301), .C1(new_n765), .C2(new_n789), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n843), .A2(G150), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G125), .C2(new_n770), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n849), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n781), .A2(G137), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G128), .A2(new_n759), .B1(new_n778), .B2(G132), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1127), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(new_n756), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n912), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n869), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n868), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n413), .B(new_n399), .C1(new_n415), .C2(new_n416), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT18), .B1(new_n417), .B2(new_n402), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1144), .B2(new_n401), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT38), .B1(new_n1145), .B2(new_n867), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT39), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n910), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1139), .B1(new_n1148), .B2(KEYINPUT100), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1138), .B1(new_n1149), .B2(new_n801), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n853), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n752), .B1(new_n370), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT120), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1123), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1122), .A2(KEYINPUT121), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT121), .B1(new_n1122), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(KEYINPUT124), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT55), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n455), .A2(new_n458), .A3(new_n463), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n461), .A2(new_n694), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1162), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n455), .A2(new_n458), .A3(new_n463), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1160), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT56), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT56), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1166), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1159), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1167), .A2(KEYINPUT56), .A3(new_n1168), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1175), .A3(KEYINPUT124), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n801), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n759), .A2(G125), .B1(G150), .B2(new_n832), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT122), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n761), .A2(G137), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n843), .A2(new_n1132), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n781), .B2(G132), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n778), .A2(G128), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT59), .Z(new_n1186));
  AOI21_X1  g0986(.A(G41), .B1(new_n827), .B2(G159), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G33), .B1(new_n770), .B2(G124), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n301), .B1(new_n268), .B2(G41), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n761), .A2(new_n338), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G41), .B(new_n330), .C1(new_n770), .C2(G283), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n843), .A2(G77), .B1(new_n827), .B2(G58), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n1004), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n217), .A2(new_n782), .B1(new_n785), .B2(new_n212), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(G107), .C2(new_n778), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT58), .Z(new_n1197));
  NAND3_X1  g0997(.A1(new_n1189), .A2(new_n1190), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n755), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n752), .B1(G50), .B2(new_n1151), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT123), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1178), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n917), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n918), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n1149), .C2(new_n905), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n887), .A2(G330), .A3(new_n897), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1177), .A2(G330), .A3(new_n897), .A4(new_n887), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n1209), .B2(new_n1208), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1202), .B1(new_n1212), .B2(new_n750), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n919), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1215), .A2(new_n1216), .B1(new_n1120), .B2(new_n1100), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n713), .B1(new_n1217), .B2(KEYINPUT57), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G375));
  AOI21_X1  g1023(.A(new_n750), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n885), .A2(new_n884), .A3(new_n801), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1151), .A2(G68), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n770), .A2(G128), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n789), .B2(new_n775), .C1(new_n301), .C2(new_n765), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G132), .B2(new_n759), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n778), .A2(G137), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n352), .B1(new_n827), .B2(G58), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n781), .A2(new_n1132), .B1(new_n761), .B2(G150), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n765), .A2(new_n339), .B1(new_n775), .B2(new_n217), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n352), .B1(new_n774), .B2(new_n769), .C1(new_n795), .C2(new_n773), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G77), .C2(new_n827), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n333), .B2(new_n798), .C1(new_n763), .C2(new_n785), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n782), .A2(new_n476), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1233), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n753), .B(new_n1226), .C1(new_n1239), .C2(new_n755), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT125), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1224), .B1(new_n1225), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1117), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1107), .A2(new_n1243), .A3(new_n962), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(G381));
  INV_X1    g1045(.A(G396), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1054), .A2(new_n1246), .A3(new_n1056), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(G387), .A2(G390), .A3(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1122), .A2(new_n1154), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1222), .A2(new_n1249), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G384), .A3(G381), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  NAND2_X1  g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1247), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n961), .A2(new_n957), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n988), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1257), .A2(new_n986), .B1(new_n973), .B2(new_n976), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n962), .B1(new_n1258), .B2(new_n744), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1256), .B1(new_n1259), .B2(new_n750), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1060), .A2(new_n1080), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1058), .A2(new_n977), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1263), .B2(new_n712), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1260), .A2(new_n1264), .A3(new_n1017), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G390), .B1(new_n991), .B2(new_n1018), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1255), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1264), .B1(new_n1260), .B2(new_n1017), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n991), .A2(new_n1018), .A3(G390), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1247), .A4(new_n1254), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n695), .A2(G213), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1222), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1120), .A2(new_n1100), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n962), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1217), .A2(KEYINPUT126), .A3(new_n962), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1249), .B1(new_n1280), .B2(new_n1213), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1272), .B1(new_n1273), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n713), .B1(new_n1243), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1107), .C1(new_n1284), .C2(new_n1243), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1242), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G384), .A2(new_n1242), .A3(new_n1286), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1282), .A2(KEYINPUT127), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1282), .B2(new_n1291), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1292), .A2(new_n1293), .A3(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1272), .A2(G2897), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1290), .B(new_n1295), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1273), .A2(new_n1281), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1272), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n1290), .B(new_n1272), .C1(new_n1273), .C2(new_n1281), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1298), .B(new_n1299), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1271), .B1(new_n1294), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1271), .B1(KEYINPUT63), .B2(new_n1301), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1303), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1249), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1273), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1291), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1271), .ZN(G402));
endmodule


