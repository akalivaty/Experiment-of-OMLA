//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT33), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(new_n206), .B2(new_n205), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210));
  AND2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(KEYINPUT23), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n212), .A2(new_n219), .A3(KEYINPUT23), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n210), .B(new_n213), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT25), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(KEYINPUT64), .A3(new_n217), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n219), .B1(new_n212), .B2(KEYINPUT23), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n232), .A3(new_n213), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n211), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n216), .B2(new_n217), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n231), .B2(new_n230), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .A3(KEYINPUT25), .A4(new_n229), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n224), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT27), .B1(new_n224), .B2(KEYINPUT66), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n227), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT27), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G183gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n224), .A2(KEYINPUT27), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n224), .A2(KEYINPUT27), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(G190gat), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n240), .B(new_n244), .C1(new_n253), .C2(new_n242), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n212), .A2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n256), .A2(KEYINPUT26), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n211), .B1(new_n256), .B2(KEYINPUT26), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(G183gat), .B2(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n251), .B1(new_n249), .B2(new_n250), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n227), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT28), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n240), .B1(new_n264), .B2(new_n244), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n239), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n267));
  INV_X1    g066(.A(G134gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(G127gat), .ZN(new_n269));
  INV_X1    g068(.A(G127gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(G134gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n267), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G113gat), .B(G120gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(G134gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(G127gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT71), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n278));
  NAND4_X1  g077(.A1(new_n272), .A2(new_n274), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n269), .A2(KEYINPUT70), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n281), .B(new_n282), .C1(KEYINPUT1), .C2(new_n273), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n279), .A2(new_n286), .A3(new_n283), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n279), .B2(new_n283), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(new_n239), .C1(new_n260), .C2(new_n265), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G227gat), .ZN(new_n295));
  INV_X1    g094(.A(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n209), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  AOI211_X1 g098(.A(KEYINPUT74), .B(new_n299), .C1(new_n289), .C2(new_n293), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT32), .B(new_n208), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT76), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n293), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n244), .B1(new_n253), .B2(new_n242), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n254), .A3(new_n259), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n292), .B1(new_n307), .B2(new_n239), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n297), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n209), .A3(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n312), .A2(KEYINPUT76), .A3(KEYINPUT32), .A4(new_n208), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT34), .B1(new_n294), .B2(new_n297), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT34), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n289), .A2(new_n316), .A3(new_n299), .A4(new_n293), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT77), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n317), .A2(KEYINPUT77), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n322));
  INV_X1    g121(.A(new_n205), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n202), .B1(new_n298), .B2(new_n300), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n314), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n321), .B1(new_n314), .B2(new_n325), .ZN(new_n327));
  OR3_X1    g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT36), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT36), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G197gat), .B(G204gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT22), .ZN(new_n332));
  INV_X1    g131(.A(G211gat), .ZN(new_n333));
  INV_X1    g132(.A(G218gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT78), .ZN(new_n339));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT79), .B(KEYINPUT29), .Z(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n266), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n307), .B2(new_n239), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n266), .A2(new_n341), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n307), .B2(new_n239), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n338), .B(new_n346), .C1(new_n347), .C2(new_n341), .ZN(new_n348));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  NAND4_X1  g150(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT30), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n345), .B2(new_n348), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n345), .A2(new_n348), .A3(new_n351), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT81), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n345), .A2(new_n348), .A3(new_n360), .A4(new_n351), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n354), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT2), .ZN(new_n366));
  INV_X1    g165(.A(G148gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(G141gat), .ZN(new_n368));
  INV_X1    g167(.A(G141gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(G148gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G155gat), .ZN(new_n372));
  INV_X1    g171(.A(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n365), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT82), .B1(new_n374), .B2(new_n365), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT83), .B1(new_n367), .B2(G141gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n369), .A3(G148gat), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n378), .B(new_n380), .C1(new_n369), .C2(G148gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n365), .B1(new_n374), .B2(KEYINPUT2), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n364), .B1(new_n288), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n279), .A2(new_n283), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n374), .A2(new_n365), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n365), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n391), .A2(new_n371), .B1(new_n381), .B2(new_n382), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n384), .A2(KEYINPUT3), .B1(new_n283), .B2(new_n279), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n398), .A3(new_n383), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n396), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n399), .A3(new_n284), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n395), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n279), .A2(new_n377), .A3(new_n383), .A4(new_n283), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT84), .B1(new_n408), .B2(KEYINPUT4), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n386), .A2(new_n392), .A3(new_n410), .A4(new_n364), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT4), .B1(new_n288), .B2(new_n384), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n407), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n284), .A2(new_n384), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n408), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n401), .B1(new_n416), .B2(new_n396), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n404), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n364), .B1(new_n292), .B2(new_n392), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n409), .A2(new_n411), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n400), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(KEYINPUT85), .A3(new_n417), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n403), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NOR2_X1   g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  INV_X1    g230(.A(new_n403), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n414), .A2(new_n404), .A3(new_n418), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT85), .B1(new_n422), .B2(new_n417), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n428), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n430), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n363), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT31), .B(G50gat), .ZN(new_n441));
  INV_X1    g240(.A(G106gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n338), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n399), .A2(new_n342), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT86), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n339), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT3), .B1(new_n338), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(G228gat), .B(G233gat), .C1(new_n454), .C2(new_n392), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G22gat), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n338), .A2(new_n342), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n384), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g259(.A(new_n338), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n447), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n460), .A2(new_n462), .B1(G228gat), .B2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n455), .B1(new_n449), .B2(new_n451), .ZN(new_n466));
  OAI21_X1  g265(.A(G22gat), .B1(new_n466), .B2(new_n463), .ZN(new_n467));
  INV_X1    g266(.A(G78gat), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n444), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n465), .A2(new_n467), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G78gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n443), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n440), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n330), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n358), .A2(new_n361), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n346), .B1(new_n347), .B2(new_n341), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n343), .A2(new_n344), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(new_n339), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT38), .B1(new_n483), .B2(KEYINPUT37), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n351), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n355), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n424), .B2(new_n428), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n424), .B2(new_n428), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n435), .A2(KEYINPUT87), .A3(new_n436), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n493), .A3(new_n430), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n488), .A2(new_n493), .A3(new_n496), .A4(new_n430), .ZN(new_n497));
  INV_X1    g296(.A(new_n487), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n485), .B1(new_n345), .B2(new_n348), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT38), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n471), .A2(new_n475), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n385), .A2(new_n406), .A3(new_n393), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n396), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(KEYINPUT39), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n504), .B(KEYINPUT39), .C1(new_n396), .C2(new_n416), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n428), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT40), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n508), .A2(new_n490), .A3(new_n492), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n354), .A2(new_n356), .A3(new_n362), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n501), .A2(new_n511), .A3(KEYINPUT89), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT89), .B1(new_n501), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n478), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n326), .A2(new_n327), .A3(new_n502), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n440), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n314), .A2(new_n325), .ZN(new_n518));
  INV_X1    g317(.A(new_n321), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n314), .A2(new_n321), .A3(new_n325), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n476), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n493), .A2(new_n430), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n363), .A3(new_n515), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n514), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(G1gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n530), .B2(G1gat), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT93), .A3(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(new_n531), .A3(new_n536), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n542), .B(new_n543), .C1(G29gat), .C2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  OAI221_X1 g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .C1(new_n539), .C2(KEYINPUT15), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT91), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT14), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n541), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G43gat), .B(G50gat), .Z(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(new_n540), .A3(new_n550), .A4(new_n544), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n552), .A2(new_n556), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI211_X1 g361(.A(KEYINPUT92), .B(KEYINPUT17), .C1(new_n552), .C2(new_n556), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n538), .B(new_n558), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n535), .A2(new_n537), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n560), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n527), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT90), .B(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT11), .B(G169gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT12), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT94), .B1(new_n557), .B2(new_n538), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n567), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n566), .A2(KEYINPUT94), .A3(new_n560), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n565), .B(KEYINPUT13), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n569), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n564), .A2(KEYINPUT18), .A3(new_n565), .A4(new_n567), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n582), .A2(new_n581), .B1(new_n568), .B2(new_n569), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n588), .B(new_n585), .C1(new_n570), .C2(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n526), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n438), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n593), .A2(G57gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(G57gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT9), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G71gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n468), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT96), .B(G57gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n594), .B1(new_n602), .B2(G64gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(KEYINPUT9), .B2(new_n599), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT20), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n566), .B1(KEYINPUT21), .B2(new_n606), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n614), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(G99gat), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT8), .B1(new_n630), .B2(new_n442), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G99gat), .B(G106gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT7), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n629), .A3(new_n631), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n633), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n641), .A2(new_n560), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n562), .A2(new_n563), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n558), .A2(new_n640), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n625), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n623), .B1(new_n646), .B2(KEYINPUT99), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n643), .A2(new_n644), .ZN(new_n648));
  INV_X1    g447(.A(new_n642), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n624), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n645), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n605), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n603), .A2(new_n604), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n637), .A2(new_n657), .A3(new_n639), .A4(new_n601), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n606), .A3(KEYINPUT100), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT10), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n655), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n655), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(new_n666), .A3(new_n661), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT101), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n667), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n618), .A2(new_n654), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n591), .A2(new_n592), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT102), .B(G1gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  AND3_X1   g479(.A1(new_n591), .A2(new_n510), .A3(new_n677), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n532), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  AND2_X1   g485(.A1(new_n591), .A2(new_n677), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n330), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n326), .A2(new_n327), .ZN(new_n690));
  INV_X1    g489(.A(new_n677), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n591), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(G1326gat));
  NAND2_X1  g493(.A1(new_n687), .A2(new_n502), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  AND2_X1   g496(.A1(new_n526), .A2(new_n654), .ZN(new_n698));
  INV_X1    g497(.A(new_n618), .ZN(new_n699));
  INV_X1    g498(.A(new_n590), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(new_n700), .A3(new_n676), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n545), .A3(new_n592), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n328), .B(new_n329), .C1(new_n476), .C2(new_n440), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n501), .A2(new_n511), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT89), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n501), .A2(new_n511), .A3(KEYINPUT89), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n517), .B2(new_n525), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT35), .B1(new_n522), .B2(new_n439), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n523), .A2(new_n363), .A3(new_n515), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n516), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n715), .A3(KEYINPUT103), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n654), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n517), .A2(new_n525), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT44), .B(new_n654), .C1(new_n710), .C2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n701), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n438), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n724), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n702), .A2(new_n546), .A3(new_n510), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n723), .B2(new_n363), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(G43gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n702), .A2(new_n731), .A3(new_n690), .ZN(new_n732));
  INV_X1    g531(.A(new_n330), .ZN(new_n733));
  OAI21_X1  g532(.A(G43gat), .B1(new_n723), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1330gat));
  NAND4_X1  g536(.A1(new_n720), .A2(new_n502), .A3(new_n701), .A4(new_n722), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G50gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n476), .A2(G50gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n698), .A2(new_n701), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n740), .B1(new_n739), .B2(new_n742), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT104), .B1(new_n738), .B2(G50gat), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n745), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n746), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n743), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1331gat));
  AND3_X1   g551(.A1(new_n713), .A2(new_n715), .A3(KEYINPUT103), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT103), .B1(new_n713), .B2(new_n715), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n514), .ZN(new_n756));
  INV_X1    g555(.A(new_n676), .ZN(new_n757));
  NOR4_X1   g556(.A1(new_n618), .A2(new_n590), .A3(new_n654), .A4(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n592), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(new_n602), .Z(G1332gat));
  INV_X1    g560(.A(KEYINPUT49), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n759), .B(new_n510), .C1(new_n762), .C2(new_n593), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n593), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(new_n759), .ZN(new_n767));
  OAI21_X1  g566(.A(G71gat), .B1(new_n767), .B2(new_n733), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n759), .A2(new_n597), .A3(new_n690), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g570(.A1(new_n759), .A2(new_n502), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n626), .A2(new_n628), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n699), .A2(new_n590), .A3(new_n757), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n720), .A2(new_n722), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(new_n438), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n699), .A2(new_n590), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n654), .B(new_n778), .C1(new_n710), .C2(new_n717), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT107), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  INV_X1    g581(.A(new_n654), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n755), .B2(new_n514), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT51), .A4(new_n778), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n757), .A2(new_n774), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n592), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n777), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n363), .A2(G92gat), .A3(new_n757), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n720), .A2(new_n510), .A3(new_n722), .A4(new_n775), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n796), .B2(G92gat), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  INV_X1    g598(.A(new_n782), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n779), .A2(new_n780), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n794), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(G92gat), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT109), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n795), .A2(new_n797), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n802), .A2(new_n803), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n799), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n776), .B2(new_n733), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n690), .A2(new_n630), .A3(new_n676), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n788), .B2(new_n812), .ZN(G1338gat));
  OR2_X1    g612(.A1(new_n776), .A2(new_n476), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n476), .A2(G106gat), .A3(new_n757), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n787), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n800), .A2(new_n801), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n814), .A2(G106gat), .B1(new_n820), .B2(new_n818), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n817), .A2(new_n819), .B1(new_n821), .B2(new_n816), .ZN(G1339gat));
  OAI21_X1  g621(.A(new_n672), .B1(new_n665), .B2(KEYINPUT54), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n665), .A2(KEYINPUT54), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n662), .A2(new_n655), .A3(new_n664), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n662), .A2(new_n664), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n666), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(KEYINPUT110), .A3(KEYINPUT54), .A4(new_n665), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n823), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT55), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n590), .A3(new_n675), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT111), .B1(new_n831), .B2(KEYINPUT55), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n827), .A2(new_n830), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n823), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n586), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n581), .A2(new_n582), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n565), .B1(new_n564), .B2(new_n567), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n840), .A2(new_n576), .B1(new_n843), .B2(new_n575), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n676), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT113), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n838), .A2(new_n834), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n848), .B(new_n845), .C1(new_n849), .C2(new_n833), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n783), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n844), .A2(new_n832), .A3(new_n654), .A4(new_n675), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n853), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n834), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(KEYINPUT112), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n699), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n691), .A2(new_n590), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n863));
  INV_X1    g662(.A(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n845), .B1(new_n849), .B2(new_n833), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n654), .B1(new_n865), .B2(KEYINPUT113), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n858), .B1(new_n866), .B2(new_n850), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n863), .B(new_n864), .C1(new_n867), .C2(new_n699), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n363), .A3(new_n592), .A4(new_n516), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n700), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n757), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g673(.A1(new_n870), .A2(new_n618), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT115), .B(G127gat), .Z(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1342gat));
  INV_X1    g676(.A(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n654), .B1(new_n878), .B2(new_n268), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n330), .A2(new_n438), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n363), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n831), .A2(KEYINPUT55), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n845), .B1(new_n833), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n783), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n854), .A2(new_n887), .A3(new_n857), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(KEYINPUT116), .A3(new_n618), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n864), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT116), .B1(new_n888), .B2(new_n618), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n502), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n862), .A2(new_n868), .A3(new_n894), .A4(new_n502), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n895), .A3(new_n590), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT58), .B1(new_n896), .B2(G141gat), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n862), .A2(new_n868), .A3(new_n502), .A4(new_n883), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n510), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n590), .A2(new_n369), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT118), .Z(new_n904));
  OAI21_X1  g703(.A(new_n897), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n896), .A2(KEYINPUT117), .A3(G141gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT117), .B1(new_n896), .B2(G141gat), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n898), .A2(new_n510), .A3(new_n904), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1344gat));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n862), .A2(new_n868), .A3(new_n502), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n855), .A2(new_n856), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n699), .B1(new_n887), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n894), .B(new_n502), .C1(new_n916), .C2(new_n861), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n884), .A2(new_n757), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n912), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n893), .A2(new_n895), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n757), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(KEYINPUT59), .A3(new_n367), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n676), .A2(new_n367), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n921), .A2(new_n924), .B1(new_n902), .B2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n922), .B2(new_n618), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n699), .A2(new_n372), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n902), .B2(new_n928), .ZN(G1346gat));
  NOR3_X1   g728(.A1(new_n922), .A2(new_n373), .A3(new_n783), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n900), .A2(new_n654), .A3(new_n901), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n373), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n592), .A2(new_n363), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n862), .A2(new_n868), .A3(new_n516), .A4(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n700), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(new_n214), .ZN(G1348gat));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n757), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(new_n215), .ZN(G1349gat));
  NOR2_X1   g737(.A1(new_n934), .A2(new_n618), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n261), .A2(new_n262), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n934), .B2(new_n618), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(KEYINPUT121), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT60), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n939), .A2(new_n947), .A3(new_n941), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n944), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n944), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(G1350gat));
  OAI22_X1  g750(.A1(new_n934), .A2(new_n783), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(G1351gat));
  XNOR2_X1  g753(.A(KEYINPUT123), .B(G197gat), .ZN(new_n955));
  INV_X1    g754(.A(new_n933), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n330), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n918), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n958), .B2(new_n700), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n330), .A2(new_n476), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n869), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n700), .A2(new_n955), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n914), .A2(new_n676), .A3(new_n917), .A4(new_n957), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(KEYINPUT125), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n966), .B1(KEYINPUT125), .B2(new_n965), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n869), .A2(new_n964), .A3(new_n676), .A4(new_n960), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(KEYINPUT62), .ZN(new_n970));
  XOR2_X1   g769(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n967), .A2(new_n972), .ZN(G1353gat));
  NAND4_X1  g772(.A1(new_n914), .A2(new_n699), .A3(new_n917), .A4(new_n957), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G211gat), .ZN(new_n975));
  NOR2_X1   g774(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n974), .B(G211gat), .C1(KEYINPUT126), .C2(KEYINPUT63), .ZN(new_n978));
  NAND2_X1  g777(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n961), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n981), .A2(new_n333), .A3(new_n699), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n958), .B2(new_n783), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n334), .A3(new_n654), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


