//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT65), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n476), .A3(G137), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n475), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n465), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n472), .C2(G112), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n472), .A2(new_n476), .A3(G138), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n472), .A2(new_n476), .A3(KEYINPUT4), .A4(G138), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n476), .A2(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n490), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n501), .A2(new_n503), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT66), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(new_n516), .A3(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(G88), .B1(new_n520), .B2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  INV_X1    g101(.A(new_n518), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n525), .B1(new_n526), .B2(new_n527), .C1(new_n532), .C2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(new_n518), .A2(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n519), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n513), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(new_n518), .A2(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n519), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n513), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n518), .A2(G91), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n508), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n514), .A2(new_n516), .A3(G53), .A4(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n560), .B2(KEYINPUT68), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NOR3_X1   g137(.A1(new_n560), .A2(KEYINPUT68), .A3(KEYINPUT9), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n555), .B(new_n559), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(G299));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n567));
  XNOR2_X1  g142(.A(G171), .B(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G301));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n513), .B1(new_n508), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT71), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n518), .A2(G87), .B1(new_n520), .B2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT72), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n501), .A2(new_n503), .A3(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n518), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n518), .A2(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n519), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n513), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  XOR2_X1   g163(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n527), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n508), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n518), .A2(G92), .A3(new_n589), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT73), .B1(new_n599), .B2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  MUX2_X1   g176(.A(KEYINPUT73), .B(new_n600), .S(new_n601), .Z(G284));
  MUX2_X1   g177(.A(KEYINPUT73), .B(new_n600), .S(new_n601), .Z(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n564), .B(KEYINPUT69), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n599), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n481), .A2(G123), .ZN(new_n614));
  OAI221_X1 g189(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n472), .C2(G111), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n484), .A2(G135), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT76), .B(G2096), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n620));
  NOR3_X1   g195(.A1(new_n463), .A2(new_n461), .A3(G2105), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT13), .B(G2100), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT15), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2435), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n630), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n638), .A2(G14), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT78), .Z(new_n646));
  XOR2_X1   g221(.A(new_n644), .B(KEYINPUT17), .Z(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n644), .A3(new_n640), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n642), .A3(new_n640), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  INV_X1    g245(.A(G1981), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(G229));
  NAND2_X1  g249(.A1(new_n599), .A2(G16), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G4), .B2(G16), .ZN(new_n676));
  INV_X1    g251(.A(G1348), .ZN(new_n677));
  INV_X1    g252(.A(G2078), .ZN(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NOR2_X1   g254(.A1(G164), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G27), .B2(new_n679), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n676), .A2(new_n677), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G5), .A2(G16), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G171), .B2(G16), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n605), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g261(.A1(new_n685), .A2(KEYINPUT23), .A3(G20), .ZN(new_n687));
  AOI21_X1  g262(.A(KEYINPUT23), .B1(new_n685), .B2(G20), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(G1956), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(G1956), .ZN(new_n691));
  OAI221_X1 g266(.A(new_n682), .B1(G1961), .B2(new_n684), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(G29), .A2(G35), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G162), .B2(G29), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(G2090), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n676), .A2(new_n677), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n692), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n681), .A2(new_n678), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G29), .A2(G33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n484), .A2(G139), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(new_n472), .C2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n702), .B1(new_n707), .B2(new_n679), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n712));
  NOR2_X1   g287(.A1(KEYINPUT24), .A2(G34), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(G160), .A2(G29), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n712), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2084), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n696), .A2(G2090), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n699), .A2(new_n701), .A3(new_n711), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G286), .A2(new_n685), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(KEYINPUT84), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(G1966), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G28), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(new_n679), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n684), .A2(G1961), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT87), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n617), .A2(new_n679), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT85), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n735), .A2(new_n736), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n708), .A2(new_n709), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n481), .A2(G129), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n484), .A2(G141), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND4_X1  g322(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G29), .B2(G32), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT27), .B(G1996), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT83), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n742), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n723), .A2(new_n741), .A3(new_n756), .ZN(new_n757));
  OAI221_X1 g332(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n472), .C2(G107), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT79), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n481), .A2(G119), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n484), .A2(G131), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G25), .B(new_n762), .S(G29), .Z(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT35), .B(G1991), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n685), .A2(G24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n587), .B2(new_n685), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1986), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT34), .ZN(new_n770));
  INV_X1    g345(.A(G288), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G23), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT33), .B(G1976), .Z(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n685), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n685), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(G1971), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(G1971), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n772), .B(new_n774), .C1(G16), .C2(G23), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n776), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT32), .B(G1981), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n782), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n783), .B1(new_n782), .B2(new_n787), .ZN(new_n789));
  AOI211_X1 g364(.A(KEYINPUT81), .B(new_n770), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n770), .A2(KEYINPUT81), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n770), .A2(KEYINPUT81), .ZN(new_n792));
  AND4_X1   g367(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n769), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(KEYINPUT36), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(new_n769), .C1(new_n790), .C2(new_n793), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n685), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n548), .B2(new_n685), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1341), .Z(new_n801));
  NOR3_X1   g376(.A1(new_n735), .A2(new_n738), .A3(new_n740), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT88), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n757), .A2(new_n798), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n751), .A2(new_n753), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n679), .A2(G26), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n481), .A2(G128), .ZN(new_n808));
  OAI221_X1 g383(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n472), .C2(G116), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n484), .A2(G140), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(new_n679), .ZN(new_n813));
  MUX2_X1   g388(.A(new_n807), .B(new_n813), .S(KEYINPUT28), .Z(new_n814));
  INV_X1    g389(.A(G2067), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n804), .A2(new_n806), .A3(new_n817), .ZN(G311));
  AND3_X1   g393(.A1(new_n757), .A2(new_n798), .A3(new_n803), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n819), .A2(new_n805), .A3(new_n816), .A4(new_n801), .ZN(G150));
  NAND2_X1  g395(.A1(new_n518), .A2(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n519), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n513), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  AOI21_X1  g404(.A(new_n547), .B1(KEYINPUT91), .B2(new_n826), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT91), .B2(new_n826), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(new_n832), .A3(new_n547), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n598), .A2(new_n608), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n829), .B1(new_n839), .B2(G860), .ZN(G145));
  XOR2_X1   g415(.A(new_n762), .B(new_n622), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n484), .A2(G142), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT95), .Z(new_n843));
  OAI221_X1 g418(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n472), .C2(G118), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n481), .A2(G130), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n841), .A2(new_n846), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT96), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(G160), .B(KEYINPUT92), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n486), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n617), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT96), .ZN(new_n856));
  OR2_X1    g431(.A1(G102), .A2(G2105), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(new_n496), .A3(G2104), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n462), .A2(new_n464), .A3(new_n492), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT93), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT93), .B1(new_n858), .B2(new_n859), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n490), .B(new_n491), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n811), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n749), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(new_n707), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n707), .B(new_n866), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n855), .A2(new_n856), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n856), .A2(new_n867), .A3(new_n869), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n853), .A3(new_n854), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g450(.A1(new_n827), .A2(G868), .ZN(new_n876));
  XNOR2_X1  g451(.A(G303), .B(new_n587), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G305), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n771), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n878), .B(G288), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n883), .A2(KEYINPUT98), .A3(KEYINPUT42), .ZN(new_n884));
  OAI22_X1  g459(.A1(new_n882), .A2(new_n884), .B1(new_n880), .B2(new_n881), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(KEYINPUT99), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n834), .B(new_n610), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n605), .A2(new_n599), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n598), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n887), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT97), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n887), .B2(new_n890), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n885), .A2(KEYINPUT99), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n886), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n885), .A2(new_n899), .A3(KEYINPUT99), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n876), .B1(new_n904), .B2(G868), .ZN(G295));
  AOI21_X1  g480(.A(new_n876), .B1(new_n904), .B2(G868), .ZN(G331));
  NOR2_X1   g481(.A1(new_n568), .A2(G286), .ZN(new_n907));
  AND2_X1   g482(.A1(G286), .A2(G171), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n834), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n833), .B(new_n831), .C1(new_n907), .C2(new_n908), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n892), .A2(new_n894), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n890), .A3(new_n911), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT100), .A3(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(KEYINPUT100), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n883), .A2(KEYINPUT101), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT101), .A4(new_n883), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n871), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n890), .A2(KEYINPUT102), .A3(new_n891), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n912), .B(new_n924), .C1(new_n913), .C2(KEYINPUT102), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n879), .B1(new_n925), .B2(new_n915), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(KEYINPUT103), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n918), .B2(new_n879), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(KEYINPUT103), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n923), .B1(new_n930), .B2(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n922), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  MUX2_X1   g509(.A(new_n931), .B(new_n934), .S(KEYINPUT44), .Z(G397));
  XOR2_X1   g510(.A(KEYINPUT104), .B(G1384), .Z(new_n936));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n862), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n474), .A2(G40), .A3(new_n478), .A4(new_n477), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n940), .A2(G1996), .A3(new_n748), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n811), .B(G2067), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT106), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(new_n748), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n940), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n945), .A2(G1996), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n942), .B(new_n943), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n762), .B(new_n764), .Z(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n940), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n940), .A2(G1986), .A3(G290), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT48), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n762), .A2(new_n764), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n812), .A2(new_n815), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n940), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n940), .A2(G1996), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT46), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n947), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n954), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n490), .A2(new_n491), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n497), .A2(KEYINPUT93), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n858), .A2(new_n859), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT93), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n939), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G8), .ZN(new_n972));
  NAND2_X1  g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n578), .A2(new_n579), .A3(new_n671), .A4(new_n580), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n973), .A2(KEYINPUT49), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT49), .B1(new_n973), .B2(new_n974), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n572), .A2(G1976), .A3(new_n573), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n971), .A2(G8), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n982), .A3(KEYINPUT52), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n498), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n862), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n939), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1971), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n938), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(G2090), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n862), .A2(new_n999), .A3(new_n989), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n988), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n987), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n979), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT108), .B(G1976), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G288), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1004), .A2(KEYINPUT109), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n971), .A2(new_n1005), .A3(G8), .A4(new_n978), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1007), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n984), .A2(new_n1003), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n862), .A2(new_n989), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n498), .A2(new_n999), .A3(new_n989), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1016), .A2(new_n939), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  AOI21_X1  g594(.A(G2090), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n938), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1017), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1020), .A2(new_n1023), .B1(new_n995), .B2(new_n994), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n986), .B1(new_n1024), .B2(new_n988), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1014), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n939), .B(new_n1027), .C1(new_n970), .C2(KEYINPUT45), .ZN(new_n1028));
  INV_X1    g603(.A(G1966), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT112), .B(G2084), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n939), .A3(new_n1000), .A4(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n997), .A2(KEYINPUT113), .A3(new_n1000), .A4(new_n1032), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1030), .A2(new_n1035), .A3(new_n1039), .A4(new_n1036), .ZN(new_n1040));
  AND2_X1   g615(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1042), .A2(G8), .A3(G286), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n1037), .B2(G8), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(G168), .A3(new_n1040), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1026), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT62), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n997), .A2(new_n1000), .ZN(new_n1053));
  INV_X1    g628(.A(G1961), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n938), .B1(new_n1015), .B2(new_n991), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2078), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1027), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(KEYINPUT122), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT122), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n994), .A2(G2078), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(KEYINPUT53), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G301), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1043), .C2(new_n1046), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1049), .A2(new_n1052), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n563), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1070), .A2(new_n561), .B1(G651), .B2(new_n558), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(KEYINPUT57), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(KEYINPUT57), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1071), .A2(new_n555), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n564), .A2(new_n1072), .A3(KEYINPUT57), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1956), .B1(new_n1021), .B2(new_n1017), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n992), .A2(new_n939), .A3(new_n993), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1077), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(new_n1080), .C1(new_n1018), .C2(G1956), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT61), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1087), .B(KEYINPUT61), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1015), .A2(new_n938), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1053), .A2(new_n677), .B1(new_n815), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g666(.A(KEYINPUT119), .B(new_n599), .C1(new_n1091), .C2(KEYINPUT60), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1053), .A2(new_n677), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n815), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n598), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1092), .A2(new_n1097), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1082), .A2(new_n1084), .A3(KEYINPUT61), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(KEYINPUT116), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n971), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1996), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n992), .A2(new_n1106), .A3(new_n993), .A4(new_n939), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT117), .B1(new_n1108), .B2(new_n548), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1111), .B(new_n547), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1103), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1103), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1109), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1089), .A2(new_n1100), .A3(new_n1101), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1082), .B1(new_n598), .B2(new_n1091), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1084), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1057), .B1(new_n994), .B2(G2078), .ZN(new_n1123));
  OAI211_X1 g698(.A(G301), .B(new_n1123), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n937), .B1(KEYINPUT123), .B2(new_n939), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n993), .A3(new_n1058), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(new_n1123), .A3(new_n1055), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(KEYINPUT54), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1124), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1129), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1128), .A2(new_n568), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1066), .B2(G301), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1136));
  AOI22_X1  g711(.A1(new_n1132), .A2(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1047), .A2(new_n1026), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1122), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1037), .A2(G8), .A3(G168), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1014), .A2(new_n1025), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n984), .A2(new_n1003), .A3(new_n1013), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT63), .B1(new_n987), .B2(new_n1002), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(new_n1142), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  AND4_X1   g721(.A1(new_n987), .A2(new_n984), .A3(new_n1002), .A4(new_n1013), .ZN(new_n1147));
  OR3_X1    g722(.A1(new_n977), .A2(G1976), .A3(G288), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT110), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1148), .A2(new_n1149), .A3(new_n974), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1148), .B2(new_n974), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n972), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1146), .A2(new_n1147), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1069), .A2(new_n1139), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n940), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n587), .B(G1986), .Z(new_n1156));
  AOI21_X1  g731(.A(new_n951), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1154), .A2(KEYINPUT126), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT126), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n963), .B1(new_n1158), .B2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g735(.A1(G401), .A2(G227), .ZN(new_n1162));
  AND2_X1   g736(.A1(new_n874), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g737(.A(G229), .ZN(new_n1164));
  NAND4_X1  g738(.A1(new_n931), .A2(new_n1163), .A3(G319), .A4(new_n1164), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


