

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752;

  NOR2_X1 U369 ( .A1(n630), .A2(n373), .ZN(n631) );
  OR2_X1 U370 ( .A1(n573), .A2(n531), .ZN(n579) );
  XNOR2_X1 U371 ( .A(n528), .B(n527), .ZN(n543) );
  XNOR2_X2 U372 ( .A(n599), .B(n512), .ZN(n610) );
  XNOR2_X2 U373 ( .A(n387), .B(KEYINPUT45), .ZN(n734) );
  NAND2_X1 U374 ( .A1(n346), .A2(n533), .ZN(n697) );
  NAND2_X1 U375 ( .A1(n385), .A2(n626), .ZN(n368) );
  AND2_X1 U376 ( .A1(n579), .A2(n580), .ZN(n391) );
  NAND2_X1 U377 ( .A1(n396), .A2(KEYINPUT66), .ZN(n395) );
  XNOR2_X1 U378 ( .A(n363), .B(n362), .ZN(n596) );
  OR2_X1 U379 ( .A1(n624), .A2(n577), .ZN(n363) );
  XNOR2_X1 U380 ( .A(n555), .B(n554), .ZN(n637) );
  AND2_X1 U381 ( .A1(n717), .A2(n412), .ZN(n411) );
  NAND2_X1 U382 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U383 ( .A(n702), .B(n360), .ZN(n564) );
  INV_X2 U384 ( .A(n692), .ZN(n346) );
  AND2_X1 U385 ( .A1(n652), .A2(n507), .ZN(n403) );
  XOR2_X1 U386 ( .A(n645), .B(KEYINPUT59), .Z(n646) );
  XNOR2_X1 U387 ( .A(n384), .B(n383), .ZN(n490) );
  XNOR2_X1 U388 ( .A(n446), .B(G119), .ZN(n384) );
  NOR2_X1 U389 ( .A1(n632), .A2(n631), .ZN(n347) );
  NOR2_X1 U390 ( .A1(n632), .A2(n631), .ZN(n349) );
  NAND2_X1 U391 ( .A1(n397), .A2(n395), .ZN(n348) );
  NOR2_X1 U392 ( .A1(n632), .A2(n631), .ZN(n350) );
  NAND2_X1 U393 ( .A1(n397), .A2(n395), .ZN(n650) );
  NOR2_X1 U394 ( .A1(n632), .A2(n631), .ZN(n651) );
  XNOR2_X2 U395 ( .A(n351), .B(G469), .ZN(n529) );
  NOR2_X1 U396 ( .A1(n663), .A2(G902), .ZN(n351) );
  XNOR2_X2 U397 ( .A(n629), .B(n628), .ZN(n632) );
  BUF_X1 U398 ( .A(n347), .Z(n662) );
  NAND2_X1 U399 ( .A1(n543), .A2(n698), .ZN(n573) );
  OR2_X1 U400 ( .A1(n652), .A2(n419), .ZN(n404) );
  XNOR2_X1 U401 ( .A(n652), .B(n653), .ZN(n654) );
  XNOR2_X2 U402 ( .A(n481), .B(n433), .ZN(n394) );
  XNOR2_X2 U403 ( .A(n392), .B(n687), .ZN(n481) );
  NAND2_X1 U404 ( .A1(n382), .A2(n381), .ZN(n598) );
  XNOR2_X1 U405 ( .A(n375), .B(n374), .ZN(n445) );
  XNOR2_X1 U406 ( .A(G146), .B(KEYINPUT98), .ZN(n374) );
  XNOR2_X1 U407 ( .A(n376), .B(KEYINPUT5), .ZN(n375) );
  NAND2_X1 U408 ( .A1(n464), .A2(G210), .ZN(n376) );
  XNOR2_X1 U409 ( .A(n425), .B(n424), .ZN(n477) );
  XOR2_X1 U410 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n425) );
  AND2_X1 U411 ( .A1(n748), .A2(n377), .ZN(n464) );
  INV_X1 U412 ( .A(G237), .ZN(n377) );
  XOR2_X1 U413 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n463) );
  XNOR2_X1 U414 ( .A(KEYINPUT4), .B(G131), .ZN(n433) );
  NAND2_X1 U415 ( .A1(n504), .A2(KEYINPUT2), .ZN(n372) );
  NAND2_X1 U416 ( .A1(n371), .A2(n734), .ZN(n370) );
  NOR2_X1 U417 ( .A1(n368), .A2(n627), .ZN(n371) );
  NAND2_X1 U418 ( .A1(n420), .A2(n627), .ZN(n419) );
  INV_X1 U419 ( .A(n507), .ZN(n420) );
  XNOR2_X1 U420 ( .A(n569), .B(n568), .ZN(n717) );
  INV_X1 U421 ( .A(G472), .ZN(n380) );
  XNOR2_X1 U422 ( .A(G113), .B(KEYINPUT3), .ZN(n383) );
  XNOR2_X1 U423 ( .A(n416), .B(G137), .ZN(n434) );
  INV_X1 U424 ( .A(G140), .ZN(n416) );
  XNOR2_X1 U425 ( .A(n415), .B(KEYINPUT83), .ZN(n414) );
  INV_X1 U426 ( .A(KEYINPUT24), .ZN(n415) );
  NAND2_X1 U427 ( .A1(n477), .A2(G221), .ZN(n417) );
  XNOR2_X1 U428 ( .A(G122), .B(G116), .ZN(n482) );
  INV_X1 U429 ( .A(G104), .ZN(n439) );
  XNOR2_X1 U430 ( .A(KEYINPUT90), .B(G110), .ZN(n440) );
  NOR2_X1 U431 ( .A1(G902), .A2(G237), .ZN(n450) );
  INV_X1 U432 ( .A(n588), .ZN(n389) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U434 ( .A(n448), .B(n447), .ZN(n639) );
  XNOR2_X1 U435 ( .A(G137), .B(G116), .ZN(n444) );
  XNOR2_X1 U436 ( .A(G131), .B(G140), .ZN(n462) );
  XOR2_X1 U437 ( .A(G122), .B(G104), .Z(n461) );
  XNOR2_X1 U438 ( .A(KEYINPUT76), .B(KEYINPUT17), .ZN(n495) );
  XNOR2_X1 U439 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n494) );
  NOR2_X1 U440 ( .A1(n712), .A2(n713), .ZN(n589) );
  AND2_X1 U441 ( .A1(n526), .A2(n570), .ZN(n412) );
  NAND2_X1 U442 ( .A1(n551), .A2(n410), .ZN(n409) );
  INV_X1 U443 ( .A(n570), .ZN(n410) );
  NAND2_X1 U444 ( .A1(n353), .A2(n379), .ZN(n704) );
  XNOR2_X1 U445 ( .A(n573), .B(KEYINPUT107), .ZN(n401) );
  NOR2_X1 U446 ( .A1(n399), .A2(n346), .ZN(n398) );
  NOR2_X1 U447 ( .A1(n702), .A2(n574), .ZN(n399) );
  XNOR2_X1 U448 ( .A(n443), .B(n369), .ZN(n378) );
  INV_X1 U449 ( .A(KEYINPUT97), .ZN(n369) );
  XOR2_X1 U450 ( .A(KEYINPUT62), .B(n639), .Z(n640) );
  INV_X1 U451 ( .A(n747), .ZN(n367) );
  XNOR2_X1 U452 ( .A(n490), .B(n489), .ZN(n493) );
  XNOR2_X1 U453 ( .A(n417), .B(n413), .ZN(n426) );
  XNOR2_X1 U454 ( .A(n434), .B(n414), .ZN(n413) );
  NOR2_X1 U455 ( .A1(n748), .A2(G952), .ZN(n668) );
  INV_X1 U456 ( .A(n630), .ZN(n690) );
  INV_X1 U457 ( .A(G134), .ZN(n687) );
  INV_X1 U458 ( .A(KEYINPUT40), .ZN(n362) );
  XOR2_X1 U459 ( .A(n422), .B(n354), .Z(n352) );
  XNOR2_X1 U460 ( .A(G902), .B(KEYINPUT15), .ZN(n627) );
  NOR2_X1 U461 ( .A1(n698), .A2(n697), .ZN(n353) );
  XOR2_X1 U462 ( .A(G119), .B(G128), .Z(n354) );
  NOR2_X1 U463 ( .A1(n546), .A2(n545), .ZN(n355) );
  NOR2_X1 U464 ( .A1(n576), .A2(KEYINPUT44), .ZN(n356) );
  OR2_X1 U465 ( .A1(n418), .A2(n510), .ZN(n357) );
  AND2_X1 U466 ( .A1(n702), .A2(n574), .ZN(n358) );
  AND2_X1 U467 ( .A1(n404), .A2(n421), .ZN(n359) );
  XOR2_X1 U468 ( .A(n530), .B(KEYINPUT6), .Z(n360) );
  XNOR2_X1 U469 ( .A(n731), .B(n503), .ZN(n652) );
  XNOR2_X1 U470 ( .A(n493), .B(n492), .ZN(n731) );
  INV_X1 U471 ( .A(KEYINPUT2), .ZN(n373) );
  XNOR2_X2 U472 ( .A(n361), .B(KEYINPUT10), .ZN(n743) );
  XNOR2_X1 U473 ( .A(n361), .B(n392), .ZN(n497) );
  XNOR2_X2 U474 ( .A(G146), .B(G125), .ZN(n361) );
  INV_X1 U475 ( .A(n596), .ZN(n382) );
  XNOR2_X1 U476 ( .A(n562), .B(n561), .ZN(n624) );
  XNOR2_X2 U477 ( .A(n364), .B(n430), .ZN(n692) );
  NAND2_X1 U478 ( .A1(n633), .A2(n485), .ZN(n364) );
  XNOR2_X1 U479 ( .A(n365), .B(n426), .ZN(n633) );
  XNOR2_X1 U480 ( .A(n423), .B(n352), .ZN(n365) );
  NAND2_X1 U481 ( .A1(n734), .A2(n366), .ZN(n630) );
  INV_X1 U482 ( .A(n368), .ZN(n366) );
  XNOR2_X1 U483 ( .A(n368), .B(n367), .ZN(n749) );
  NAND2_X1 U484 ( .A1(n370), .A2(n372), .ZN(n629) );
  NAND2_X2 U485 ( .A1(n402), .A2(n404), .ZN(n599) );
  NAND2_X1 U486 ( .A1(n389), .A2(n356), .ZN(n388) );
  XNOR2_X1 U487 ( .A(n550), .B(n549), .ZN(n575) );
  NAND2_X1 U488 ( .A1(n590), .A2(n379), .ZN(n591) );
  NOR2_X1 U489 ( .A1(n702), .A2(n510), .ZN(n452) );
  NAND2_X1 U490 ( .A1(n378), .A2(n702), .ZN(n521) );
  INV_X1 U491 ( .A(n702), .ZN(n379) );
  XNOR2_X2 U492 ( .A(n449), .B(n380), .ZN(n702) );
  INV_X1 U493 ( .A(n752), .ZN(n381) );
  XNOR2_X1 U494 ( .A(n386), .B(n623), .ZN(n385) );
  NAND2_X1 U495 ( .A1(n622), .A2(n621), .ZN(n386) );
  NAND2_X1 U496 ( .A1(n390), .A2(n388), .ZN(n387) );
  XNOR2_X1 U497 ( .A(n586), .B(KEYINPUT87), .ZN(n390) );
  NAND2_X1 U498 ( .A1(n581), .A2(n391), .ZN(n583) );
  XNOR2_X1 U499 ( .A(n744), .B(n442), .ZN(n663) );
  XNOR2_X2 U500 ( .A(G143), .B(G128), .ZN(n392) );
  NAND2_X1 U501 ( .A1(n359), .A2(n393), .ZN(n509) );
  INV_X1 U502 ( .A(n403), .ZN(n393) );
  XNOR2_X2 U503 ( .A(n394), .B(n435), .ZN(n744) );
  XNOR2_X1 U504 ( .A(n394), .B(n490), .ZN(n447) );
  INV_X1 U505 ( .A(n401), .ZN(n396) );
  AND2_X2 U506 ( .A1(n400), .A2(n398), .ZN(n397) );
  NAND2_X1 U507 ( .A1(n401), .A2(n358), .ZN(n400) );
  NOR2_X1 U508 ( .A1(n403), .A2(n357), .ZN(n402) );
  INV_X1 U509 ( .A(n526), .ZN(n551) );
  NAND2_X1 U510 ( .A1(n407), .A2(n405), .ZN(n572) );
  NAND2_X1 U511 ( .A1(n406), .A2(n410), .ZN(n405) );
  INV_X1 U512 ( .A(n717), .ZN(n406) );
  NOR2_X1 U513 ( .A1(n411), .A2(n408), .ZN(n407) );
  NAND2_X1 U514 ( .A1(n409), .A2(n571), .ZN(n408) );
  INV_X1 U515 ( .A(n421), .ZN(n418) );
  NAND2_X1 U516 ( .A1(n507), .A2(n504), .ZN(n421) );
  INV_X1 U517 ( .A(n510), .ZN(n511) );
  XNOR2_X1 U518 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n519) );
  INV_X1 U519 ( .A(KEYINPUT66), .ZN(n574) );
  INV_X1 U520 ( .A(n704), .ZN(n552) );
  INV_X1 U521 ( .A(n658), .ZN(n659) );
  XNOR2_X1 U522 ( .A(n743), .B(KEYINPUT95), .ZN(n423) );
  XOR2_X1 U523 ( .A(KEYINPUT23), .B(G110), .Z(n422) );
  INV_X2 U524 ( .A(G953), .ZN(n748) );
  NAND2_X1 U525 ( .A1(G234), .A2(n748), .ZN(n424) );
  INV_X1 U526 ( .A(G902), .ZN(n485) );
  NAND2_X1 U527 ( .A1(n627), .A2(G234), .ZN(n428) );
  XNOR2_X1 U528 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n428), .B(n427), .ZN(n431) );
  NAND2_X1 U530 ( .A1(G217), .A2(n431), .ZN(n429) );
  XNOR2_X1 U531 ( .A(KEYINPUT25), .B(n429), .ZN(n430) );
  AND2_X1 U532 ( .A1(n431), .A2(G221), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n432), .B(KEYINPUT21), .ZN(n533) );
  INV_X1 U534 ( .A(n533), .ZN(n693) );
  XNOR2_X1 U535 ( .A(n434), .B(KEYINPUT94), .ZN(n435) );
  NAND2_X1 U536 ( .A1(n748), .A2(G227), .ZN(n436) );
  XNOR2_X1 U537 ( .A(n436), .B(G146), .ZN(n438) );
  XNOR2_X1 U538 ( .A(G101), .B(G107), .ZN(n437) );
  XNOR2_X1 U539 ( .A(n438), .B(n437), .ZN(n441) );
  XNOR2_X1 U540 ( .A(n440), .B(n439), .ZN(n489) );
  XNOR2_X1 U541 ( .A(n441), .B(n489), .ZN(n442) );
  NOR2_X1 U542 ( .A1(n697), .A2(n529), .ZN(n443) );
  XNOR2_X1 U543 ( .A(n445), .B(n444), .ZN(n448) );
  XNOR2_X2 U544 ( .A(G101), .B(KEYINPUT68), .ZN(n446) );
  NAND2_X1 U545 ( .A1(n639), .A2(n485), .ZN(n449) );
  XNOR2_X1 U546 ( .A(n450), .B(KEYINPUT73), .ZN(n505) );
  AND2_X1 U547 ( .A1(n505), .A2(G214), .ZN(n510) );
  XOR2_X1 U548 ( .A(KEYINPUT113), .B(KEYINPUT30), .Z(n451) );
  XNOR2_X1 U549 ( .A(n452), .B(n451), .ZN(n458) );
  XNOR2_X1 U550 ( .A(n453), .B(KEYINPUT14), .ZN(n455) );
  NAND2_X1 U551 ( .A1(G952), .A2(n455), .ZN(n723) );
  NOR2_X1 U552 ( .A1(G953), .A2(n723), .ZN(n515) );
  AND2_X1 U553 ( .A1(G953), .A2(G902), .ZN(n454) );
  NAND2_X1 U554 ( .A1(n455), .A2(n454), .ZN(n513) );
  XOR2_X1 U555 ( .A(n513), .B(KEYINPUT111), .Z(n456) );
  NOR2_X1 U556 ( .A1(G900), .A2(n456), .ZN(n457) );
  OR2_X1 U557 ( .A1(n515), .A2(n457), .ZN(n532) );
  AND2_X1 U558 ( .A1(n458), .A2(n532), .ZN(n459) );
  AND2_X1 U559 ( .A1(n378), .A2(n459), .ZN(n559) );
  XNOR2_X1 U560 ( .A(G113), .B(G143), .ZN(n460) );
  XNOR2_X1 U561 ( .A(n461), .B(n460), .ZN(n468) );
  XNOR2_X1 U562 ( .A(n463), .B(n462), .ZN(n466) );
  NAND2_X1 U563 ( .A1(G214), .A2(n464), .ZN(n465) );
  XNOR2_X1 U564 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U565 ( .A(n468), .B(n467), .Z(n473) );
  XOR2_X1 U566 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n470) );
  XNOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT99), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U569 ( .A(n743), .B(n471), .Z(n472) );
  XNOR2_X1 U570 ( .A(n473), .B(n472), .ZN(n645) );
  NOR2_X1 U571 ( .A1(G902), .A2(n645), .ZN(n475) );
  XNOR2_X1 U572 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U574 ( .A(n476), .B(G475), .ZN(n557) );
  AND2_X1 U575 ( .A1(n477), .A2(G217), .ZN(n480) );
  XOR2_X1 U576 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n478) );
  XNOR2_X1 U577 ( .A(n478), .B(KEYINPUT9), .ZN(n479) );
  XNOR2_X1 U578 ( .A(n480), .B(n479), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n482), .B(G107), .ZN(n491) );
  XNOR2_X1 U580 ( .A(n481), .B(n491), .ZN(n483) );
  XNOR2_X1 U581 ( .A(n484), .B(n483), .ZN(n658) );
  NAND2_X1 U582 ( .A1(n658), .A2(n485), .ZN(n487) );
  INV_X1 U583 ( .A(G478), .ZN(n486) );
  XNOR2_X1 U584 ( .A(n487), .B(n486), .ZN(n524) );
  OR2_X1 U585 ( .A1(n557), .A2(n524), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n488), .B(KEYINPUT109), .ZN(n571) );
  XNOR2_X1 U587 ( .A(n491), .B(KEYINPUT16), .ZN(n492) );
  XNOR2_X1 U588 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n497), .B(n496), .ZN(n502) );
  XOR2_X1 U590 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n500) );
  NAND2_X1 U591 ( .A1(G224), .A2(n748), .ZN(n498) );
  XNOR2_X1 U592 ( .A(n498), .B(KEYINPUT75), .ZN(n499) );
  XNOR2_X1 U593 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U594 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U595 ( .A(n627), .ZN(n504) );
  NAND2_X1 U596 ( .A1(n505), .A2(G210), .ZN(n506) );
  XNOR2_X1 U597 ( .A(n506), .B(KEYINPUT80), .ZN(n507) );
  INV_X1 U598 ( .A(n509), .ZN(n541) );
  AND2_X1 U599 ( .A1(n571), .A2(n541), .ZN(n508) );
  NAND2_X1 U600 ( .A1(n559), .A2(n508), .ZN(n606) );
  XNOR2_X1 U601 ( .A(n606), .B(G143), .ZN(G45) );
  XNOR2_X1 U602 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n512) );
  NOR2_X1 U603 ( .A1(G898), .A2(n513), .ZN(n514) );
  OR2_X1 U604 ( .A1(n515), .A2(n514), .ZN(n517) );
  INV_X1 U605 ( .A(KEYINPUT93), .ZN(n516) );
  XNOR2_X1 U606 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X1 U607 ( .A1(n610), .A2(n518), .ZN(n520) );
  XNOR2_X2 U608 ( .A(n520), .B(n519), .ZN(n526) );
  OR2_X1 U609 ( .A1(n551), .A2(n521), .ZN(n670) );
  INV_X1 U610 ( .A(n524), .ZN(n556) );
  OR2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n577) );
  XNOR2_X1 U612 ( .A(n577), .B(KEYINPUT110), .ZN(n680) );
  NOR2_X1 U613 ( .A1(n670), .A2(n680), .ZN(n523) );
  XNOR2_X1 U614 ( .A(G104), .B(KEYINPUT115), .ZN(n522) );
  XNOR2_X1 U615 ( .A(n523), .B(n522), .ZN(G6) );
  NAND2_X1 U616 ( .A1(n557), .A2(n524), .ZN(n712) );
  NOR2_X1 U617 ( .A1(n712), .A2(n693), .ZN(n525) );
  NAND2_X1 U618 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U619 ( .A(KEYINPUT22), .ZN(n527) );
  XNOR2_X2 U620 ( .A(n529), .B(KEYINPUT1), .ZN(n698) );
  INV_X1 U621 ( .A(KEYINPUT105), .ZN(n530) );
  NAND2_X1 U622 ( .A1(n564), .A2(n346), .ZN(n531) );
  XNOR2_X1 U623 ( .A(n579), .B(G101), .ZN(G3) );
  INV_X1 U624 ( .A(n698), .ZN(n602) );
  INV_X1 U625 ( .A(n532), .ZN(n535) );
  NAND2_X1 U626 ( .A1(n692), .A2(n533), .ZN(n534) );
  NOR2_X1 U627 ( .A1(n535), .A2(n534), .ZN(n590) );
  NOR2_X1 U628 ( .A1(n680), .A2(n564), .ZN(n536) );
  NAND2_X1 U629 ( .A1(n590), .A2(n536), .ZN(n600) );
  INV_X1 U630 ( .A(n600), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n511), .A2(n537), .ZN(n538) );
  OR2_X1 U632 ( .A1(n602), .A2(n538), .ZN(n540) );
  XOR2_X1 U633 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n539) );
  XNOR2_X1 U634 ( .A(n540), .B(n539), .ZN(n542) );
  OR2_X1 U635 ( .A1(n542), .A2(n541), .ZN(n625) );
  XNOR2_X1 U636 ( .A(n625), .B(G140), .ZN(G42) );
  XNOR2_X1 U637 ( .A(n564), .B(KEYINPUT79), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n602), .A2(n692), .ZN(n544) );
  XNOR2_X1 U639 ( .A(n544), .B(KEYINPUT106), .ZN(n545) );
  NAND2_X1 U640 ( .A1(n543), .A2(n355), .ZN(n550) );
  XNOR2_X1 U641 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n548) );
  INV_X1 U642 ( .A(KEYINPUT65), .ZN(n547) );
  XNOR2_X1 U643 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n575), .B(G119), .ZN(G21) );
  INV_X1 U645 ( .A(n551), .ZN(n553) );
  INV_X1 U646 ( .A(KEYINPUT31), .ZN(n554) );
  NAND2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n674) );
  NOR2_X1 U648 ( .A1(n637), .A2(n674), .ZN(n558) );
  XOR2_X1 U649 ( .A(G116), .B(n558), .Z(G18) );
  XNOR2_X1 U650 ( .A(n509), .B(KEYINPUT38), .ZN(n710) );
  NAND2_X1 U651 ( .A1(n559), .A2(n710), .ZN(n562) );
  INV_X1 U652 ( .A(KEYINPUT70), .ZN(n560) );
  XNOR2_X1 U653 ( .A(n560), .B(KEYINPUT39), .ZN(n561) );
  XOR2_X1 U654 ( .A(G131), .B(n596), .Z(G33) );
  NOR2_X2 U655 ( .A1(n697), .A2(n698), .ZN(n563) );
  XNOR2_X1 U656 ( .A(n563), .B(KEYINPUT108), .ZN(n566) );
  INV_X1 U657 ( .A(n564), .ZN(n565) );
  NAND2_X1 U658 ( .A1(n566), .A2(n565), .ZN(n569) );
  INV_X1 U659 ( .A(KEYINPUT69), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n567), .B(KEYINPUT33), .ZN(n568) );
  XNOR2_X1 U661 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n570) );
  XNOR2_X2 U662 ( .A(n572), .B(KEYINPUT35), .ZN(n576) );
  XOR2_X1 U663 ( .A(n576), .B(G122), .Z(G24) );
  NAND2_X1 U664 ( .A1(n650), .A2(n575), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n587), .A2(KEYINPUT44), .ZN(n585) );
  NAND2_X1 U666 ( .A1(n576), .A2(KEYINPUT44), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n637), .A2(n670), .ZN(n578) );
  NAND2_X1 U668 ( .A1(n577), .A2(n674), .ZN(n604) );
  NAND2_X1 U669 ( .A1(n578), .A2(n604), .ZN(n580) );
  INV_X1 U670 ( .A(KEYINPUT88), .ZN(n582) );
  XNOR2_X1 U671 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n585), .A2(n584), .ZN(n586) );
  BUF_X1 U673 ( .A(n587), .Z(n588) );
  NAND2_X1 U674 ( .A1(n710), .A2(n511), .ZN(n713) );
  XNOR2_X1 U675 ( .A(n589), .B(KEYINPUT41), .ZN(n724) );
  XOR2_X1 U676 ( .A(KEYINPUT28), .B(KEYINPUT114), .Z(n592) );
  XNOR2_X1 U677 ( .A(n592), .B(n591), .ZN(n594) );
  INV_X1 U678 ( .A(n529), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n594), .A2(n593), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n724), .A2(n609), .ZN(n595) );
  XNOR2_X1 U681 ( .A(n595), .B(KEYINPUT42), .ZN(n752) );
  INV_X1 U682 ( .A(KEYINPUT46), .ZN(n597) );
  XNOR2_X1 U683 ( .A(n598), .B(n597), .ZN(n622) );
  NOR2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U685 ( .A(n601), .B(KEYINPUT36), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n685) );
  XNOR2_X1 U687 ( .A(n685), .B(KEYINPUT86), .ZN(n615) );
  INV_X1 U688 ( .A(n604), .ZN(n714) );
  NAND2_X1 U689 ( .A1(KEYINPUT47), .A2(n714), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n605), .B(KEYINPUT82), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U692 ( .A(n608), .B(KEYINPUT81), .ZN(n613) );
  INV_X1 U693 ( .A(n609), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n681) );
  NAND2_X1 U695 ( .A1(n681), .A2(KEYINPUT47), .ZN(n612) );
  AND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n620) );
  INV_X1 U698 ( .A(n681), .ZN(n676) );
  NOR2_X1 U699 ( .A1(KEYINPUT47), .A2(n714), .ZN(n616) );
  XNOR2_X1 U700 ( .A(KEYINPUT72), .B(n616), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n676), .A2(n617), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n618), .B(KEYINPUT71), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U704 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n623) );
  OR2_X1 U705 ( .A1(n624), .A2(n674), .ZN(n688) );
  AND2_X1 U706 ( .A1(n688), .A2(n625), .ZN(n626) );
  INV_X1 U707 ( .A(KEYINPUT64), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n662), .A2(G217), .ZN(n635) );
  INV_X1 U709 ( .A(n633), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n636), .A2(n668), .ZN(G66) );
  NOR2_X1 U712 ( .A1(n637), .A2(n680), .ZN(n638) );
  XOR2_X1 U713 ( .A(G113), .B(n638), .Z(G15) );
  NAND2_X1 U714 ( .A1(n350), .A2(G472), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n642), .A2(n668), .ZN(n644) );
  XNOR2_X1 U717 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n644), .B(n643), .ZN(G57) );
  NAND2_X1 U719 ( .A1(n349), .A2(G475), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n648), .A2(n668), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U723 ( .A(n348), .B(G110), .ZN(G12) );
  NAND2_X1 U724 ( .A1(n651), .A2(G210), .ZN(n655) );
  XOR2_X1 U725 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n653) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n656), .A2(n668), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U729 ( .A1(n662), .A2(G478), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n661), .A2(n668), .ZN(G63) );
  NAND2_X1 U732 ( .A1(n662), .A2(G469), .ZN(n667) );
  XNOR2_X1 U733 ( .A(KEYINPUT125), .B(KEYINPUT57), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT58), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n663), .B(n665), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n669) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(G54) );
  NOR2_X1 U738 ( .A1(n670), .A2(n674), .ZN(n672) );
  XNOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U741 ( .A(G107), .B(n673), .ZN(G9) );
  XOR2_X1 U742 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n678) );
  INV_X1 U743 ( .A(n674), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U746 ( .A(G128), .B(n679), .ZN(G30) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U748 ( .A(G146), .B(KEYINPUT117), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(G48) );
  XOR2_X1 U750 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n684) );
  XNOR2_X1 U751 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U752 ( .A(G125), .B(n686), .ZN(G27) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U754 ( .A(n689), .B(KEYINPUT119), .ZN(G36) );
  XOR2_X1 U755 ( .A(KEYINPUT53), .B(KEYINPUT124), .Z(n730) );
  XNOR2_X1 U756 ( .A(n690), .B(n373), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n691), .A2(G953), .ZN(n728) );
  XOR2_X1 U758 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n695) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U761 ( .A(KEYINPUT120), .B(n696), .ZN(n701) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U763 ( .A(KEYINPUT50), .B(n699), .Z(n700) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n706), .B(KEYINPUT123), .ZN(n708) );
  XOR2_X1 U768 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n707) );
  XNOR2_X1 U769 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n724), .A2(n709), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n710), .A2(n511), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n718), .A2(n406), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U777 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n724), .A2(n406), .ZN(n725) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n730), .B(n729), .ZN(G75) );
  INV_X1 U783 ( .A(G898), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(G953), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n731), .A2(n732), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n733), .B(KEYINPUT126), .ZN(n742) );
  AND2_X1 U787 ( .A1(n734), .A2(n748), .ZN(n739) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n735) );
  XOR2_X1 U789 ( .A(KEYINPUT61), .B(n735), .Z(n736) );
  NOR2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U792 ( .A(n740), .B(KEYINPUT127), .Z(n741) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n744), .B(n743), .ZN(n747) );
  XOR2_X1 U795 ( .A(G227), .B(n747), .Z(n745) );
  NAND2_X1 U796 ( .A1(G900), .A2(n745), .ZN(n746) );
  NAND2_X1 U797 ( .A1(n746), .A2(G953), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U800 ( .A(G137), .B(n752), .Z(G39) );
endmodule

