//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G229gat), .A2(G233gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT13), .Z(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(G50gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G43gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR3_X1   g016(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT15), .B(new_n215), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n212), .B2(new_n214), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(G43gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n211), .A2(G50gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT15), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  INV_X1    g027(.A(G29gat), .ZN(new_n229));
  INV_X1    g028(.A(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n216), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n224), .A2(new_n227), .A3(new_n232), .A4(new_n220), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT95), .ZN(new_n235));
  INV_X1    g034(.A(G15gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G22gat), .ZN(new_n237));
  INV_X1    g036(.A(G22gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G15gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT94), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(G15gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT94), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n235), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n241), .B2(new_n242), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n245), .A2(G1gat), .B1(new_n248), .B2(KEYINPUT16), .ZN(new_n249));
  INV_X1    g048(.A(G1gat), .ZN(new_n250));
  AOI211_X1 g049(.A(new_n235), .B(new_n250), .C1(new_n240), .C2(new_n244), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n249), .A2(G8gat), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G8gat), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT95), .B1(new_n246), .B2(new_n247), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(new_n244), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT16), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n254), .A2(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n245), .A2(G1gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n234), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(G8gat), .B1(new_n249), .B2(new_n251), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n253), .A3(new_n258), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(new_n234), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n210), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n222), .A2(KEYINPUT17), .A3(new_n233), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT96), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT96), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n222), .A2(new_n233), .A3(new_n269), .A4(KEYINPUT17), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT93), .B(KEYINPUT17), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n234), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n271), .A2(new_n262), .A3(new_n263), .A4(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n260), .A3(KEYINPUT97), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n268), .A2(new_n270), .B1(new_n234), .B2(new_n272), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT97), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n262), .A4(new_n263), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n275), .A2(new_n278), .B1(G229gat), .B2(G233gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n266), .B1(new_n279), .B2(KEYINPUT18), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n278), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n281), .A2(KEYINPUT18), .A3(new_n209), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n208), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n209), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT18), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n279), .A2(KEYINPUT18), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n266), .A4(new_n207), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n288), .A3(KEYINPUT98), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT98), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(new_n208), .C1(new_n280), .C2(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(new_n238), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  XOR2_X1   g095(.A(G141gat), .B(G148gat), .Z(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT2), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT80), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G155gat), .B(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n301), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n297), .B(new_n300), .C1(KEYINPUT80), .C2(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n296), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G211gat), .A2(G218gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(KEYINPUT75), .B2(KEYINPUT22), .ZN(new_n317));
  AND2_X1   g116(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(KEYINPUT89), .ZN(new_n323));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(KEYINPUT89), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n321), .B2(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n311), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n321), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT3), .B1(new_n329), .B2(new_n296), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n309), .A2(KEYINPUT81), .A3(new_n310), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n322), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G228gat), .A3(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G78gat), .B(G106gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(new_n213), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT88), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n328), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n328), .B2(new_n336), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n295), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n294), .A3(new_n341), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT70), .B(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT71), .ZN(new_n351));
  INV_X1    g150(.A(G113gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G120gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G127gat), .B(G134gat), .Z(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT1), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n353), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n349), .B2(G113gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G113gat), .B(G120gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT69), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT1), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n363), .B2(new_n362), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n357), .A2(new_n361), .B1(new_n355), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n309), .A2(new_n310), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n363), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n355), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n356), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n360), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n369), .B1(new_n376), .B2(new_n311), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n332), .A2(KEYINPUT3), .A3(new_n333), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n367), .A2(new_n312), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n376), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n368), .B(new_n377), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT39), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  AND2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n384), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n367), .B(new_n374), .C1(new_n360), .C2(new_n375), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n392), .B(new_n393), .C1(new_n334), .C2(new_n366), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n376), .A2(new_n332), .A3(KEYINPUT83), .A4(new_n333), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n391), .B(KEYINPUT39), .C1(new_n396), .C2(new_n384), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n390), .A2(new_n397), .A3(KEYINPUT40), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT40), .B1(new_n390), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n376), .A2(new_n332), .A3(new_n333), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n393), .B1(new_n376), .B2(new_n311), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n384), .B(new_n395), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n394), .A2(KEYINPUT84), .A3(new_n384), .A4(new_n395), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n376), .B(new_n379), .C1(new_n334), .C2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(new_n383), .A3(new_n377), .A4(new_n368), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(KEYINPUT85), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(KEYINPUT5), .A3(new_n412), .ZN(new_n415));
  INV_X1    g214(.A(new_n389), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n400), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G8gat), .B(G36gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT79), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G183gat), .ZN(new_n428));
  INV_X1    g227(.A(G190gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT24), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(new_n426), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G169gat), .ZN(new_n435));
  INV_X1    g234(.A(G176gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n435), .A2(new_n436), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n439), .A2(G169gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(new_n436), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n428), .A3(new_n429), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n432), .A2(new_n446), .A3(new_n425), .A4(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT65), .B(G176gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n442), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n440), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n434), .A2(new_n444), .B1(new_n451), .B2(new_n441), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT26), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT26), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(G169gat), .B2(G176gat), .ZN(new_n455));
  OAI221_X1 g254(.A(new_n453), .B1(new_n428), .B2(new_n429), .C1(new_n438), .C2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT27), .B(G183gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n429), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT67), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(KEYINPUT28), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n457), .B(new_n429), .C1(new_n459), .C2(KEYINPUT28), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n424), .B1(new_n464), .B2(KEYINPUT29), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT77), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT77), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(new_n424), .C1(new_n464), .C2(KEYINPUT29), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT78), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n462), .ZN(new_n471));
  INV_X1    g270(.A(new_n456), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT68), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n452), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n470), .B1(new_n477), .B2(new_n424), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n444), .A2(new_n434), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n451), .A2(new_n441), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n471), .A2(new_n475), .A3(new_n472), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n475), .B1(new_n471), .B2(new_n472), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n424), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT78), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n469), .A2(new_n329), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n464), .A2(new_n424), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n424), .B1(new_n477), .B2(KEYINPUT29), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(KEYINPUT76), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n484), .B2(new_n296), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n329), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n423), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n492), .A2(new_n493), .B1(new_n424), .B2(new_n464), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n490), .A2(KEYINPUT76), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n321), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n469), .A2(new_n329), .A3(new_n487), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n422), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(KEYINPUT30), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(new_n503), .A3(new_n500), .A4(new_n422), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n348), .B1(new_n418), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n410), .A2(KEYINPUT5), .A3(new_n412), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n412), .B1(new_n410), .B2(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n389), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n417), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n422), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n500), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(new_n423), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT38), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n469), .A2(new_n487), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT37), .B1(new_n522), .B2(new_n329), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n321), .B1(new_n491), .B2(new_n494), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n516), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n517), .B1(new_n499), .B2(new_n500), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT38), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n466), .A2(new_n468), .B1(new_n478), .B2(new_n486), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n517), .B1(new_n529), .B2(new_n321), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n329), .B1(new_n497), .B2(new_n498), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT38), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n422), .B1(new_n499), .B2(new_n500), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n532), .B(KEYINPUT90), .C1(new_n533), .C2(new_n518), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n526), .A2(new_n528), .A3(new_n501), .A4(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n507), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n513), .A2(new_n514), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n348), .B1(new_n537), .B2(new_n506), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT34), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n484), .A2(new_n366), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n376), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n544), .ZN(new_n546));
  AOI211_X1 g345(.A(KEYINPUT34), .B(new_n546), .C1(new_n541), .C2(new_n542), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G43gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT72), .ZN(new_n550));
  INV_X1    g349(.A(G71gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G99gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(new_n546), .A3(new_n542), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT33), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(KEYINPUT32), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n554), .B(KEYINPUT32), .C1(new_n555), .C2(new_n553), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n548), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT74), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT74), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n548), .A2(new_n558), .A3(new_n562), .A4(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n558), .A2(new_n559), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n539), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n548), .B1(new_n558), .B2(new_n559), .ZN(new_n570));
  AOI211_X1 g369(.A(KEYINPUT36), .B(new_n570), .C1(new_n561), .C2(new_n563), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n536), .A2(new_n538), .A3(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n564), .A2(new_n347), .A3(new_n568), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n515), .A2(new_n574), .A3(new_n505), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n570), .B1(new_n561), .B2(new_n563), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n505), .A2(new_n577), .A3(new_n578), .A4(new_n347), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n537), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n292), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT104), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(G57gat), .A2(G64gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT99), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT100), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n262), .B(new_n263), .C1(new_n594), .C2(new_n593), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT101), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT7), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(KEYINPUT101), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n613), .A2(new_n621), .A3(new_n615), .A4(new_n619), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n623), .B(new_n624), .C1(new_n591), .C2(new_n592), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n624), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n593), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT10), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n625), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n637), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n276), .A2(new_n631), .ZN(new_n646));
  INV_X1    g445(.A(new_n631), .ZN(new_n647));
  AND2_X1   g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n647), .A2(new_n234), .B1(KEYINPUT41), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G190gat), .B(G218gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n654), .A3(new_n649), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n656), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n608), .A2(new_n645), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n582), .A2(new_n583), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n400), .A2(new_n417), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n347), .B1(new_n667), .B2(new_n505), .ZN(new_n668));
  AND4_X1   g467(.A1(new_n501), .A2(new_n526), .A3(new_n528), .A4(new_n534), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n537), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n513), .A2(new_n514), .B1(new_n504), .B2(new_n502), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n572), .B1(new_n671), .B2(new_n347), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n578), .B1(new_n671), .B2(new_n574), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n537), .A2(new_n579), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n670), .A2(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n292), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n665), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT104), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n666), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n537), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AOI21_X1  g481(.A(new_n583), .B1(new_n582), .B2(new_n665), .ZN(new_n683));
  AND4_X1   g482(.A1(new_n583), .A2(new_n675), .A3(new_n676), .A4(new_n665), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n506), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n505), .B1(new_n666), .B2(new_n678), .ZN(new_n687));
  OAI22_X1  g486(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n253), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n687), .B2(new_n682), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT106), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n687), .A2(new_n253), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n687), .A2(KEYINPUT42), .A3(new_n682), .ZN(new_n693));
  INV_X1    g492(.A(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n685), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n692), .A2(new_n693), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n691), .A2(new_n697), .ZN(G1325gat));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n236), .A3(new_n577), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n572), .B1(new_n666), .B2(new_n678), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n236), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n679), .A2(new_n348), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(new_n608), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n645), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n292), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n675), .B2(new_n664), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n664), .A2(KEYINPUT107), .ZN(new_n711));
  INV_X1    g510(.A(new_n663), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n661), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n709), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n573), .B2(new_n581), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n537), .B(new_n708), .C1(new_n710), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G29gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n707), .A2(new_n713), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n515), .A2(G29gat), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n675), .A2(new_n676), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT108), .Z(G1328gat));
  AND3_X1   g525(.A1(new_n675), .A2(new_n676), .A3(new_n721), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n230), .A3(new_n506), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT46), .Z(new_n729));
  OR2_X1    g528(.A1(new_n710), .A2(new_n718), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n708), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n731), .B2(new_n505), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(new_n572), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n734), .B(new_n708), .C1(new_n710), .C2(new_n718), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n727), .A2(new_n211), .A3(new_n577), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g538(.A1(new_n727), .A2(new_n348), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n213), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n348), .A2(G50gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g543(.A(new_n675), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n608), .A2(new_n664), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n292), .A3(new_n645), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n537), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g549(.A1(new_n745), .A2(new_n505), .A3(new_n747), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  AOI21_X1  g554(.A(new_n551), .B1(new_n748), .B2(new_n734), .ZN(new_n756));
  INV_X1    g555(.A(new_n577), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(G71gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n748), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n748), .A2(new_n348), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT109), .B(G78gat), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n676), .A2(new_n705), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n645), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT110), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n730), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n617), .B1(new_n767), .B2(new_n537), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n675), .A2(new_n664), .A3(new_n764), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT51), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n675), .A2(new_n771), .A3(new_n664), .A4(new_n764), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n645), .A3(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(G85gat), .A3(new_n515), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n768), .A2(new_n774), .ZN(G1336gat));
  NOR2_X1   g574(.A1(new_n505), .A2(G92gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n770), .A2(new_n645), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n506), .B(new_n766), .C1(new_n710), .C2(new_n718), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(new_n618), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n777), .B2(KEYINPUT111), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n780), .B(new_n782), .ZN(G1337gat));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n734), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G99gat), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n757), .A2(G99gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n773), .B2(new_n786), .ZN(G1338gat));
  OAI211_X1 g586(.A(new_n348), .B(new_n766), .C1(new_n710), .C2(new_n718), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n789), .B2(KEYINPUT112), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n347), .A2(G106gat), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n770), .A2(new_n645), .A3(new_n772), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n789), .B(new_n792), .C1(KEYINPUT112), .C2(KEYINPUT53), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n633), .A2(new_n632), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT10), .B1(new_n625), .B2(new_n626), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n636), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT54), .A3(new_n634), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n642), .B1(new_n634), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n797), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808));
  INV_X1    g607(.A(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n801), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(new_n797), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n798), .A2(new_n799), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n630), .A3(new_n803), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n801), .A2(new_n814), .A3(KEYINPUT55), .A4(new_n642), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n809), .A2(new_n817), .A3(KEYINPUT55), .A4(new_n801), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n816), .A2(new_n818), .A3(new_n644), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n812), .A2(new_n289), .A3(new_n291), .A4(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n206), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n281), .A2(new_n209), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n261), .A2(new_n265), .A3(new_n210), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n288), .A2(new_n645), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n716), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n711), .A2(new_n715), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n819), .B1(new_n811), .B2(new_n807), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n288), .A2(new_n824), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n608), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n645), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n746), .A2(new_n292), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n515), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(new_n505), .A3(new_n574), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n352), .A3(new_n676), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n506), .A2(new_n757), .A3(new_n348), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n292), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  OAI21_X1  g642(.A(G120gat), .B1(new_n839), .B2(new_n832), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n835), .A2(new_n349), .A3(new_n645), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n839), .B2(new_n608), .ZN(new_n847));
  INV_X1    g646(.A(G127gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n835), .A2(new_n848), .A3(new_n705), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1342gat));
  OAI21_X1  g649(.A(G134gat), .B1(new_n839), .B2(new_n713), .ZN(new_n851));
  INV_X1    g650(.A(G134gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n852), .A3(new_n664), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n853), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT117), .B1(new_n853), .B2(KEYINPUT56), .ZN(new_n855));
  OAI221_X1 g654(.A(new_n851), .B1(KEYINPUT56), .B2(new_n853), .C1(new_n854), .C2(new_n855), .ZN(G1343gat));
  AOI21_X1  g655(.A(new_n347), .B1(new_n831), .B2(new_n833), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n572), .A2(new_n537), .A3(new_n505), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G141gat), .B1(new_n860), .B2(new_n676), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n347), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n644), .A2(new_n816), .A3(new_n818), .A4(new_n806), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n289), .A2(new_n291), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n664), .B1(new_n866), .B2(new_n825), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n828), .A2(new_n829), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n716), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n608), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n864), .B1(new_n873), .B2(new_n833), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n874), .A2(new_n875), .B1(new_n858), .B2(new_n862), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n873), .A2(new_n833), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT119), .B1(new_n877), .B2(new_n864), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n859), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n292), .A2(new_n302), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n861), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT58), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(new_n880), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n859), .B(new_n884), .C1(new_n876), .C2(new_n878), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n861), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n882), .A2(new_n886), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n860), .A2(new_n303), .A3(new_n645), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n828), .A2(new_n713), .A3(new_n829), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n608), .B1(new_n867), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n833), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n891), .B2(new_n348), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n864), .B1(new_n831), .B2(new_n833), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n859), .A2(new_n832), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G148gat), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT59), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n303), .A2(KEYINPUT59), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n879), .B2(new_n645), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n888), .B1(new_n902), .B2(new_n904), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n860), .A2(new_n298), .A3(new_n705), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n879), .A2(new_n705), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n298), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n860), .B2(new_n664), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n827), .A2(new_n299), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n879), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n910), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n859), .B(new_n914), .C1(new_n876), .C2(new_n878), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT121), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n537), .A2(new_n505), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n831), .B2(new_n833), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(new_n574), .ZN(new_n921));
  AOI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n676), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n757), .A2(new_n348), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n435), .A3(new_n292), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n922), .A2(new_n925), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n921), .B2(new_n645), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n924), .A2(new_n449), .A3(new_n832), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  NAND3_X1  g728(.A1(new_n921), .A2(new_n457), .A3(new_n705), .ZN(new_n930));
  OAI21_X1  g729(.A(G183gat), .B1(new_n924), .B2(new_n608), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n934), .B(new_n935), .Z(G1350gat));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n429), .A3(new_n716), .ZN(new_n937));
  OAI21_X1  g736(.A(G190gat), .B1(new_n924), .B2(new_n713), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(KEYINPUT61), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(KEYINPUT61), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n919), .A2(new_n734), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n857), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n676), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n572), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT123), .B1(new_n918), .B2(new_n572), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n892), .B2(new_n893), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n676), .A2(G197gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  AOI21_X1  g750(.A(G204gat), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n943), .A2(new_n645), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n948), .B2(new_n832), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1353gat));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n705), .ZN(new_n958));
  OAI21_X1  g757(.A(G211gat), .B1(new_n894), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  INV_X1    g759(.A(G211gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n961), .A3(new_n705), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1354gat));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(KEYINPUT125), .B(new_n947), .C1(new_n892), .C2(new_n893), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n664), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G218gat), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n827), .A2(G218gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n943), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n964), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n971), .ZN(new_n973));
  AOI211_X1 g772(.A(KEYINPUT126), .B(new_n973), .C1(new_n968), .C2(G218gat), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n972), .A2(new_n974), .ZN(G1355gat));
endmodule


