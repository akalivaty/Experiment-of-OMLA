//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(KEYINPUT65), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n213), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT66), .B(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n207), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n210), .B(new_n221), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G68), .Z(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n214), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT8), .A2(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT69), .B(G58), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(KEYINPUT8), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT65), .A2(G20), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT65), .A2(G20), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(G33), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n251), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n202), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n250), .B1(new_n267), .B2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n269), .B2(new_n202), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n215), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT68), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT68), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(G223), .A3(G1698), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(new_n223), .C2(new_n290), .ZN(new_n294));
  INV_X1    g0094(.A(new_n280), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n283), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n272), .B(new_n273), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n272), .A2(new_n273), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(new_n296), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n302), .A2(new_n303), .A3(new_n299), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n304), .A2(G179), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n296), .A2(G169), .B1(new_n261), .B2(new_n270), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n286), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT70), .B(G107), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n280), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G232), .A2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G238), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n320), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n281), .A2(new_n222), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n278), .B2(new_n276), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n265), .A2(new_n223), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n269), .B2(new_n223), .ZN(new_n332));
  XOR2_X1   g0132(.A(KEYINPUT8), .B(G58), .Z(new_n333));
  OR2_X1    g0133(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n257), .A2(G33), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n336), .B1(new_n223), .B2(new_n257), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n332), .B1(new_n339), .B2(new_n250), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n327), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n330), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n340), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G200), .B2(new_n327), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n328), .A2(G190), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G226), .A2(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G232), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n315), .A2(new_n316), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n295), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n279), .B1(new_n281), .B2(new_n322), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n280), .B1(new_n353), .B2(new_n354), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT13), .B1(new_n361), .B2(new_n358), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(G190), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G68), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n337), .B2(new_n223), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n250), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(KEYINPUT11), .A3(new_n250), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n371), .A2(new_n372), .B1(G68), .B2(new_n268), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n297), .B1(new_n360), .B2(new_n362), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n349), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n377), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n379), .A2(KEYINPUT72), .A3(new_n375), .A4(new_n363), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n307), .A2(new_n311), .A3(new_n348), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT78), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n254), .A2(new_n265), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n254), .B2(new_n269), .ZN(new_n385));
  XOR2_X1   g0185(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n386));
  OAI21_X1  g0186(.A(new_n217), .B1(new_n288), .B2(new_n289), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n218), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT3), .B(G33), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n285), .A2(new_n287), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n394), .A2(new_n257), .A3(KEYINPUT76), .A4(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n364), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n259), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(KEYINPUT69), .A2(G58), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT69), .A2(G58), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n211), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n404), .B2(G20), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n386), .B1(new_n397), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT74), .B1(new_n286), .B2(G33), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT74), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n284), .A3(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n410), .A3(new_n287), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT7), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G68), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n388), .B1(new_n411), .B2(new_n217), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n405), .B(KEYINPUT16), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n416), .A2(new_n250), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n385), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n410), .A2(new_n287), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n282), .A2(new_n291), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n419), .A2(KEYINPUT77), .A3(new_n408), .A4(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n408), .A2(new_n420), .A3(new_n410), .A4(new_n287), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT77), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G87), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n291), .A2(G223), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(new_n408), .A3(new_n410), .A4(new_n287), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n421), .A2(new_n424), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n295), .ZN(new_n429));
  INV_X1    g0229(.A(G190), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n279), .B1(new_n281), .B2(new_n351), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n428), .B2(new_n295), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(G200), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT17), .B1(new_n418), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n383), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n341), .B1(new_n429), .B2(new_n432), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n329), .B(new_n431), .C1(new_n428), .C2(new_n295), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT18), .B1(new_n418), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n429), .A2(G179), .A3(new_n432), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n341), .B2(new_n434), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n416), .A2(new_n250), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n387), .A2(new_n388), .B1(new_n393), .B2(new_n395), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n405), .B1(new_n447), .B2(new_n364), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n448), .B2(new_n386), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n444), .B(new_n445), .C1(new_n449), .C2(new_n385), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  INV_X1    g0252(.A(new_n385), .ZN(new_n453));
  INV_X1    g0253(.A(new_n386), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT7), .B1(new_n317), .B2(new_n217), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n393), .A2(new_n395), .ZN(new_n456));
  OAI21_X1  g0256(.A(G68), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(new_n405), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n458), .B2(new_n446), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n434), .A2(G200), .ZN(new_n460));
  AOI211_X1 g0260(.A(G190), .B(new_n431), .C1(new_n428), .C2(new_n295), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n452), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n435), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(KEYINPUT78), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n438), .A2(new_n451), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT14), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n357), .B1(new_n356), .B2(new_n359), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n361), .A2(KEYINPUT13), .A3(new_n358), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(G169), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n360), .A2(G179), .A3(new_n362), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n360), .A2(new_n362), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n467), .B1(new_n473), .B2(G169), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT73), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(G169), .B1(new_n468), .B2(new_n469), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT14), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT73), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n471), .A4(new_n470), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n375), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n382), .A2(new_n466), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n265), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n267), .A2(G33), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n251), .A2(new_n264), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n482), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n398), .A2(new_n223), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT6), .ZN(new_n490));
  AND2_X1   g0290(.A1(G97), .A2(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n487), .B(new_n489), .C1(new_n496), .C2(new_n257), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n257), .B1(new_n493), .B2(new_n495), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT79), .B1(new_n498), .B2(new_n488), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n499), .C1(new_n447), .C2(new_n319), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n486), .B1(new_n500), .B2(new_n250), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n408), .A2(new_n410), .A3(new_n291), .A4(new_n287), .ZN(new_n503));
  INV_X1    g0303(.A(G244), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n502), .A2(new_n504), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n315), .A2(new_n291), .A3(new_n316), .A4(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n315), .A2(G250), .A3(G1698), .A4(new_n316), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n295), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT81), .B1(new_n512), .B2(G41), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  INV_X1    g0314(.A(G41), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT5), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G45), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(G1), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(G41), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(KEYINPUT80), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n267), .B(G45), .C1(new_n515), .C2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND4_X1   g0324(.A1(new_n276), .A2(new_n517), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT80), .B1(new_n519), .B2(new_n520), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n516), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n295), .B1(new_n528), .B2(new_n521), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n525), .B1(new_n529), .B2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n511), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n501), .B(new_n532), .C1(new_n430), .C2(new_n531), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n319), .B1(new_n389), .B2(new_n396), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n497), .A2(new_n499), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n250), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n486), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n531), .A2(new_n341), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n511), .A2(new_n530), .A3(new_n329), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n317), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n411), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .A3(G87), .A4(new_n257), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G20), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n220), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT23), .B1(new_n318), .B2(new_n217), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n544), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g0353(.A(KEYINPUT84), .B(KEYINPUT24), .Z(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n544), .A2(new_n552), .A3(new_n554), .A4(new_n546), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n250), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n517), .A2(new_n521), .A3(new_n524), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(G264), .A3(new_n280), .ZN(new_n560));
  INV_X1    g0360(.A(G250), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n291), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G257), .B2(new_n291), .ZN(new_n563));
  INV_X1    g0363(.A(G294), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n411), .A2(new_n563), .B1(new_n284), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n295), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n528), .A2(new_n276), .A3(new_n521), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(G190), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n265), .A2(new_n494), .ZN(new_n570));
  NOR2_X1   g0370(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  INV_X1    g0374(.A(new_n485), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n572), .A2(new_n574), .B1(G107), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n560), .A2(new_n566), .A3(new_n568), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n558), .A2(new_n569), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n533), .A2(new_n541), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n264), .A2(G116), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n575), .B2(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n284), .A2(G97), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n218), .A2(new_n583), .A3(new_n219), .A4(new_n509), .ZN(new_n584));
  INV_X1    g0384(.A(G116), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n249), .A2(new_n214), .B1(G20), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n341), .B1(new_n582), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n419), .A2(G257), .A3(new_n291), .A4(new_n408), .ZN(new_n593));
  OAI21_X1  g0393(.A(G303), .B1(new_n288), .B2(new_n289), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(G264), .A2(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n408), .A2(new_n410), .A3(new_n287), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT83), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n280), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n559), .A2(new_n280), .ZN(new_n601));
  INV_X1    g0401(.A(G270), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n568), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(KEYINPUT21), .B(new_n592), .C1(new_n600), .C2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n419), .A2(new_n598), .A3(new_n408), .A4(new_n596), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n597), .A2(KEYINPUT83), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n593), .A2(new_n605), .A3(new_n594), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n295), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n525), .B1(new_n529), .B2(G270), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n582), .A2(new_n591), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .A4(G179), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n609), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT21), .B1(new_n613), .B2(new_n592), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n558), .A2(new_n576), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n577), .A2(G179), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n341), .B2(new_n577), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n613), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n297), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n613), .A2(new_n430), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n622), .A2(new_n610), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n338), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n264), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n419), .A2(G68), .A3(new_n257), .A4(new_n408), .ZN(new_n627));
  OR2_X1    g0427(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n628));
  NAND2_X1  g0428(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n354), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n543), .A2(new_n482), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n630), .A2(new_n220), .B1(new_n631), .B2(new_n318), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n218), .A2(G33), .A3(G97), .A4(new_n219), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n628), .A3(new_n629), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n627), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n635), .B2(new_n250), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n575), .A2(new_n625), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(G238), .A2(G1698), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n504), .B2(G1698), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n287), .A3(new_n408), .A4(new_n410), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n280), .B1(new_n641), .B2(new_n547), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n561), .B1(new_n518), .B2(G1), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n267), .A2(new_n274), .A3(G45), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n280), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(G169), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n504), .A2(G1698), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(G238), .B2(G1698), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n547), .B1(new_n411), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n295), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(G179), .A3(new_n645), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n638), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n575), .A2(G87), .ZN(new_n655));
  OAI21_X1  g0455(.A(G200), .B1(new_n642), .B2(new_n646), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n651), .A2(G190), .A3(new_n645), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n636), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n624), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n481), .A2(new_n580), .A3(new_n620), .A4(new_n660), .ZN(G372));
  NAND2_X1  g0461(.A1(new_n475), .A2(new_n479), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n374), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n376), .A2(new_n377), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n343), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n438), .A3(new_n465), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n451), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n310), .B1(new_n667), .B2(new_n307), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n511), .A2(new_n329), .A3(new_n530), .ZN(new_n669));
  AOI21_X1  g0469(.A(G169), .B1(new_n511), .B2(new_n530), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n501), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT86), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n341), .B1(new_n651), .B2(new_n645), .ZN(new_n673));
  AOI211_X1 g0473(.A(new_n329), .B(new_n646), .C1(new_n650), .C2(new_n295), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n647), .A2(new_n652), .A3(KEYINPUT86), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n485), .A2(new_n543), .ZN(new_n678));
  AOI211_X1 g0478(.A(new_n626), .B(new_n678), .C1(new_n635), .C2(new_n250), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n656), .A2(new_n657), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n677), .A2(new_n638), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n671), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n673), .A2(new_n674), .A3(new_n672), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT86), .B1(new_n647), .B2(new_n652), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n638), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT26), .B1(new_n541), .B2(new_n659), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT87), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n683), .A2(new_n687), .A3(KEYINPUT87), .A4(new_n686), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n658), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n615), .B2(new_n619), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n580), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n481), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n668), .A2(new_n696), .ZN(G369));
  NAND2_X1  g0497(.A1(new_n257), .A2(new_n263), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G343), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n610), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n615), .B(new_n704), .Z(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n624), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n616), .A2(new_n618), .A3(new_n702), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n558), .A2(new_n576), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n579), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n709), .B1(new_n619), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n615), .A2(new_n703), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n709), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n208), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n267), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n318), .A2(G116), .A3(new_n631), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n721), .A2(new_n722), .B1(new_n213), .B2(new_n720), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  NAND3_X1  g0524(.A1(new_n608), .A2(new_n609), .A3(G179), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT88), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT88), .A4(G179), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n642), .A2(new_n646), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n511), .A2(new_n567), .A3(new_n530), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n731), .B1(new_n727), .B2(new_n728), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT30), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n730), .A2(G179), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n531), .A2(new_n613), .A3(new_n577), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n735), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n740), .B2(new_n703), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n734), .B(new_n731), .C1(new_n727), .C2(new_n728), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT31), .B(new_n703), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT89), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n703), .B1(new_n742), .B2(new_n743), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT89), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n744), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n620), .A2(new_n660), .A3(new_n580), .A4(new_n702), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n688), .A2(new_n689), .B1(new_n580), .B2(new_n693), .ZN(new_n755));
  AOI211_X1 g0555(.A(KEYINPUT29), .B(new_n703), .C1(new_n755), .C2(new_n691), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT29), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT90), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n501), .A2(new_n670), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n680), .A2(new_n679), .B1(new_n638), .B2(new_n653), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n759), .A2(new_n760), .A3(new_n682), .A4(new_n540), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n686), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n682), .B1(new_n671), .B2(new_n681), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT26), .B1(new_n692), .B2(new_n541), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(KEYINPUT90), .A3(new_n686), .A4(new_n761), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(new_n766), .A3(new_n694), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n757), .B1(new_n767), .B2(new_n702), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n724), .B1(new_n771), .B2(G1), .ZN(G364));
  NOR2_X1   g0572(.A1(new_n220), .A2(new_n262), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G45), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n721), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n707), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n706), .A2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n214), .B1(G20), .B2(new_n341), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n411), .A2(new_n208), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n518), .B2(new_n213), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n518), .B2(new_n247), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n317), .A2(new_n719), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n788), .A2(G355), .B1(new_n585), .B2(new_n719), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n784), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n297), .A2(G179), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n792), .A2(new_n217), .A3(new_n430), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G303), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n317), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n257), .A2(new_n329), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G190), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  INV_X1    g0600(.A(G329), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G179), .A2(G200), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n220), .A2(new_n430), .A3(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n430), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n796), .B(new_n804), .C1(G322), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n257), .A2(new_n792), .A3(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT91), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT91), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n797), .A2(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G190), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT33), .B(G317), .Z(new_n818));
  OAI221_X1 g0618(.A(new_n808), .B1(new_n809), .B2(new_n814), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n815), .A2(new_n430), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n802), .A2(G190), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n220), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n820), .A2(G326), .B1(G294), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT92), .Z(new_n824));
  INV_X1    g0624(.A(new_n822), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n482), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n317), .B(new_n826), .C1(G87), .C2(new_n793), .ZN(new_n827));
  INV_X1    g0627(.A(new_n799), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G77), .A2(new_n828), .B1(new_n807), .B2(new_n253), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G50), .A2(new_n820), .B1(new_n816), .B2(G68), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n814), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G107), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n803), .A2(new_n399), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT32), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n819), .A2(new_n824), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n790), .B1(new_n837), .B2(new_n782), .ZN(new_n838));
  INV_X1    g0638(.A(new_n781), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n706), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n775), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n778), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT93), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  AOI21_X1  g0645(.A(new_n703), .B1(new_n755), .B2(new_n691), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n703), .A2(new_n345), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT95), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n344), .A2(new_n848), .A3(new_n703), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT95), .B1(new_n343), .B2(new_n702), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n348), .A2(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n703), .B(new_n851), .C1(new_n755), .C2(new_n691), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n754), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n841), .B1(new_n856), .B2(new_n754), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n851), .A2(new_n779), .ZN(new_n860));
  INV_X1    g0660(.A(new_n782), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n780), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n841), .B1(G77), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n816), .B(KEYINPUT94), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G283), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n814), .A2(new_n543), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n799), .A2(new_n585), .B1(new_n800), .B2(new_n803), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(G294), .B2(new_n807), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n317), .B1(new_n794), .B2(new_n494), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n826), .B(new_n871), .C1(G303), .C2(new_n820), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n866), .A2(new_n868), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G159), .A2(new_n828), .B1(new_n807), .B2(G143), .ZN(new_n874));
  INV_X1    g0674(.A(G150), .ZN(new_n875));
  INV_X1    g0675(.A(G137), .ZN(new_n876));
  INV_X1    g0676(.A(new_n820), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n874), .B1(new_n817), .B2(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT34), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n814), .A2(new_n364), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n253), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n545), .B1(new_n825), .B2(new_n883), .C1(new_n794), .C2(new_n202), .ZN(new_n884));
  INV_X1    g0684(.A(new_n803), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n884), .B1(G132), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n878), .A2(new_n879), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n863), .B1(new_n889), .B2(new_n782), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n858), .A2(new_n859), .B1(new_n860), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  NOR2_X1   g0692(.A1(new_n773), .A2(new_n267), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n459), .A2(new_n444), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n418), .A2(new_n435), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n701), .B1(new_n449), .B2(new_n385), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n894), .A2(new_n895), .A3(new_n896), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n463), .A2(new_n442), .A3(new_n450), .A4(new_n464), .ZN(new_n902));
  INV_X1    g0702(.A(new_n896), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n414), .A2(new_n415), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n454), .B1(new_n906), .B2(new_n405), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n453), .B1(new_n907), .B2(new_n446), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n701), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n444), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n895), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n466), .A2(new_n910), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n905), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n375), .A2(new_n702), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n664), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n663), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n381), .A2(new_n479), .A3(new_n475), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n916), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n851), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n749), .A2(new_n752), .A3(new_n744), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT40), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT98), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT40), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  AOI221_X4 g0728(.A(new_n928), .B1(new_n900), .B2(new_n913), .C1(new_n466), .C2(new_n910), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n466), .A2(new_n910), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n913), .A2(new_n900), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n927), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n921), .B2(new_n922), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n924), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(G330), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n481), .A2(new_n922), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(G330), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT99), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n937), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(KEYINPUT99), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n930), .A2(new_n931), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n928), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n930), .A2(KEYINPUT38), .A3(new_n931), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(KEYINPUT39), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n929), .B2(new_n905), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n663), .A2(new_n703), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n946), .A2(new_n947), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n918), .A2(new_n920), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n695), .A2(new_n702), .A3(new_n852), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n343), .A2(new_n703), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n953), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n451), .A2(new_n701), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n481), .B1(new_n756), .B2(new_n768), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n668), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n893), .B1(new_n944), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n944), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n496), .B(KEYINPUT96), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n968), .A2(G116), .A3(new_n215), .A4(new_n220), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT36), .Z(new_n972));
  NAND3_X1  g0772(.A1(new_n213), .A2(G77), .A3(new_n403), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n974), .A2(KEYINPUT97), .B1(new_n202), .B2(G68), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(KEYINPUT97), .B2(new_n974), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(G1), .A3(new_n262), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n966), .A2(new_n972), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT100), .ZN(G367));
  OAI221_X1 g0779(.A(new_n783), .B1(new_n208), .B2(new_n338), .C1(new_n240), .C2(new_n785), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n841), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n681), .B1(new_n679), .B2(new_n702), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n679), .A2(new_n702), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n686), .B2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n807), .A2(G303), .B1(G317), .B2(new_n885), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n482), .B2(new_n811), .C1(new_n809), .C2(new_n799), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n793), .A2(G116), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT106), .Z(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n411), .B1(new_n825), .B2(new_n319), .C1(new_n987), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G311), .B2(new_n820), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n986), .B(new_n994), .C1(G294), .C2(new_n865), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n794), .A2(new_n883), .B1(new_n876), .B2(new_n803), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT107), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n290), .B1(new_n825), .B2(new_n364), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G50), .B2(new_n828), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n807), .A2(G150), .B1(G77), .B2(new_n810), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1000), .C1(new_n1001), .C2(new_n877), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n997), .B(new_n1002), .C1(G159), .C2(new_n865), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n981), .B1(new_n839), .B2(new_n984), .C1(new_n1005), .C2(new_n861), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n774), .A2(G1), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n533), .B(new_n541), .C1(new_n501), .C2(new_n702), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n671), .A2(new_n703), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n717), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT104), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT104), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n717), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n717), .A2(new_n1010), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT44), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1012), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n714), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1017), .A2(new_n1019), .A3(new_n715), .A4(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n712), .B(new_n716), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n707), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n771), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n720), .B(KEYINPUT41), .Z(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1007), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT101), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n541), .B1(new_n1008), .B2(new_n619), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n702), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n712), .A2(new_n1010), .A3(new_n716), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT42), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1031), .B(new_n1033), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT101), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT102), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n984), .B(KEYINPUT43), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1010), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n715), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT102), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1038), .A2(new_n1050), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(KEYINPUT103), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1043), .A2(new_n1051), .A3(new_n1046), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1049), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT103), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1052), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1006), .B1(new_n1030), .B2(new_n1058), .ZN(G387));
  OAI22_X1  g0859(.A1(new_n794), .A2(new_n564), .B1(new_n809), .B2(new_n825), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n820), .A2(G322), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G303), .A2(new_n828), .B1(new_n807), .B2(G317), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n864), .C2(new_n800), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n885), .A2(G326), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n411), .C1(new_n585), .C2(new_n811), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT110), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n799), .A2(new_n364), .B1(new_n875), .B2(new_n803), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n816), .A2(new_n254), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n822), .A2(new_n625), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n411), .B1(new_n793), .B2(G77), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1072), .B(new_n1076), .C1(G50), .C2(new_n807), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n820), .A2(KEYINPUT109), .A3(G159), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n832), .A2(G97), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT109), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n877), .B2(new_n399), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n861), .B1(new_n1071), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n712), .A2(new_n839), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n237), .A2(new_n518), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n788), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1085), .A2(new_n785), .B1(new_n722), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n333), .A2(new_n202), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT50), .Z(new_n1089));
  AOI21_X1  g0889(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n722), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1087), .A2(new_n1091), .B1(new_n494), .B2(new_n719), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n841), .B1(new_n1092), .B2(new_n784), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT108), .ZN(new_n1094));
  OR3_X1    g0894(.A1(new_n1083), .A2(new_n1084), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1007), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n770), .A2(new_n1026), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n770), .A2(KEYINPUT111), .A3(new_n1026), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n720), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT111), .B1(new_n770), .B2(new_n1026), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1095), .B1(new_n1096), .B2(new_n1026), .C1(new_n1100), .C2(new_n1101), .ZN(G393));
  NAND3_X1  g0902(.A1(new_n1022), .A2(new_n1007), .A3(new_n1023), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n783), .B1(new_n482), .B2(new_n208), .C1(new_n244), .C2(new_n785), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n841), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n799), .A2(new_n564), .B1(new_n825), .B2(new_n585), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n865), .B2(G303), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT112), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n820), .A2(G317), .B1(new_n807), .B2(G311), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT52), .Z(new_n1110));
  OAI21_X1  g0910(.A(new_n317), .B1(new_n794), .B2(new_n809), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G322), .B2(new_n885), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n833), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n820), .A2(G150), .B1(new_n807), .B2(G159), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT51), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n865), .A2(G50), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n825), .A2(new_n223), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n411), .B(new_n1117), .C1(G68), .C2(new_n793), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n828), .A2(new_n333), .B1(G143), .B2(new_n885), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n868), .A2(new_n1116), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1108), .A2(new_n1113), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1105), .B1(new_n1121), .B2(new_n782), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n839), .B2(new_n1010), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n720), .B1(new_n1024), .B2(new_n1098), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1097), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1103), .B(new_n1123), .C1(new_n1124), .C2(new_n1125), .ZN(G390));
  NAND3_X1  g0926(.A1(new_n962), .A2(new_n938), .A3(new_n668), .ZN(new_n1127));
  INV_X1    g0927(.A(G330), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n851), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n954), .B1(new_n753), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n922), .A2(new_n954), .A3(new_n1129), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n958), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n767), .A2(new_n702), .A3(new_n852), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n957), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n954), .B1(new_n922), .B2(new_n1129), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n753), .A2(new_n954), .A3(new_n1129), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1127), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n954), .B1(new_n854), .B2(new_n956), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n951), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1140), .A2(new_n1141), .B1(new_n948), .B2(new_n950), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n954), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1133), .B2(new_n957), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1144), .A2(new_n951), .A3(new_n915), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1131), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1134), .A2(new_n954), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n915), .A2(new_n951), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n901), .A2(new_n904), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n928), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT39), .B1(new_n947), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n929), .A2(new_n932), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(KEYINPUT39), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n951), .B1(new_n958), .B2(new_n954), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1137), .B(new_n1149), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1139), .A2(new_n1146), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n720), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT113), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1139), .B(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n956), .B1(new_n846), .B2(new_n852), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1141), .B1(new_n1161), .B2(new_n1143), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n948), .A2(new_n950), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1162), .A2(new_n1163), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1131), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1158), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1156), .B(new_n1007), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n841), .B1(new_n254), .B2(new_n862), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n793), .A2(G150), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT53), .Z(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n290), .C1(new_n399), .C2(new_n825), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G128), .B2(new_n820), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n811), .A2(new_n202), .ZN(new_n1175));
  INV_X1    g0975(.A(G132), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1176), .A2(new_n806), .B1(new_n799), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(G125), .C2(new_n885), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1174), .B(new_n1179), .C1(new_n864), .C2(new_n876), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n864), .A2(new_n319), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n799), .A2(new_n482), .B1(new_n564), .B2(new_n803), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G116), .B2(new_n807), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n317), .B1(new_n794), .B2(new_n543), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1117), .B(new_n1184), .C1(G283), .C2(new_n820), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n882), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1180), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1170), .B1(new_n1187), .B2(new_n782), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1154), .B2(new_n780), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1169), .A2(KEYINPUT114), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT114), .B1(new_n1169), .B2(new_n1189), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT115), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1169), .A2(new_n1189), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT114), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT115), .B1(new_n1197), .B2(new_n1190), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1168), .B1(new_n1194), .B2(new_n1198), .ZN(G378));
  INV_X1    g0999(.A(new_n701), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n271), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n307), .A2(new_n311), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n307), .B2(new_n311), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OR3_X1    g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n936), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n961), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1210), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n935), .A2(G330), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n923), .A2(KEYINPUT98), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n953), .A2(new_n1216), .A3(new_n927), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1128), .B(new_n1210), .C1(new_n1217), .C2(new_n924), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1213), .B1(new_n935), .B2(G330), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n961), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1215), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1007), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n411), .A2(new_n515), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n794), .A2(new_n223), .B1(new_n364), .B2(new_n825), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n820), .C2(G116), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n482), .B2(new_n817), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n810), .A2(new_n253), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n809), .B2(new_n803), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n494), .A2(new_n806), .B1(new_n799), .B2(new_n338), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT116), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT58), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1223), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n817), .A2(new_n1176), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n794), .A2(new_n1177), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT117), .Z(new_n1236));
  AOI22_X1  g1036(.A1(new_n807), .A2(G128), .B1(G150), .B2(new_n822), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n876), .C2(new_n799), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1234), .B(new_n1238), .C1(G125), .C2(new_n820), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n810), .A2(G159), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G33), .B(G41), .C1(new_n885), .C2(G124), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1232), .B(new_n1233), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1231), .A2(KEYINPUT58), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n782), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT118), .Z(new_n1249));
  OAI21_X1  g1049(.A(new_n841), .B1(G50), .B2(new_n862), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT119), .Z(new_n1251));
  NOR2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1210), .A2(new_n779), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1222), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n720), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1127), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1215), .A2(new_n1220), .B1(new_n1157), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1258), .B2(KEYINPUT57), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1166), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1221), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1255), .B1(new_n1259), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(G375));
  NAND3_X1  g1067(.A1(new_n1132), .A2(new_n1127), .A3(new_n1138), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1160), .A2(new_n1029), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1096), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT123), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1143), .A2(new_n779), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT120), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n865), .A2(G116), .B1(new_n318), .B2(new_n828), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT121), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n832), .A2(G77), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n806), .A2(new_n809), .B1(new_n795), .B2(new_n803), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n317), .B(new_n1074), .C1(new_n794), .C2(new_n482), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1279), .B(new_n1280), .C1(G294), .C2(new_n820), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n411), .B1(new_n793), .B2(G159), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n202), .B2(new_n825), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n807), .A2(G137), .B1(G128), .B2(new_n885), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1227), .C1(new_n875), .C2(new_n799), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1284), .B(new_n1286), .C1(G132), .C2(new_n820), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n864), .B2(new_n1177), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT122), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n782), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1292));
  OAI221_X1 g1092(.A(new_n841), .B1(G68), .B2(new_n862), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1273), .A2(new_n1293), .ZN(new_n1294));
  OR3_X1    g1094(.A1(new_n1270), .A2(new_n1271), .A3(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1271), .B1(new_n1270), .B2(new_n1294), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1269), .A2(new_n1297), .ZN(G381));
  INV_X1    g1098(.A(G390), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n891), .ZN(new_n1300));
  OR2_X1    g1100(.A1(G393), .A2(G396), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(G381), .A2(new_n1300), .A3(new_n1301), .A4(G387), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1197), .A2(new_n1190), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1167), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1266), .A3(new_n1304), .ZN(G407));
  INV_X1    g1105(.A(G213), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G343), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1266), .A2(new_n1304), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G407), .A2(G213), .A3(new_n1308), .ZN(G409));
  NOR2_X1   g1109(.A1(new_n1139), .A2(new_n1256), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1132), .A2(new_n1127), .A3(KEYINPUT60), .A4(new_n1138), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1268), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1310), .A2(KEYINPUT125), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1297), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n891), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1316), .A2(new_n1297), .A3(G384), .A4(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1307), .A2(G2897), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1266), .A2(G378), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1221), .A2(new_n1029), .A3(new_n1262), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT124), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI22_X1  g1131(.A1(new_n1221), .A2(new_n1007), .B1(new_n1253), .B2(new_n1252), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1221), .A2(KEYINPUT124), .A3(new_n1262), .A4(new_n1029), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1304), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1328), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1307), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1307), .B1(new_n1328), .B2(new_n1335), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1321), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  OAI211_X1 g1144(.A(G390), .B(new_n1006), .C1(new_n1030), .C2(new_n1058), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(KEYINPUT126), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(G393), .B(G396), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G387), .A2(new_n1299), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1345), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT126), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1349), .A2(new_n1347), .A3(new_n1352), .A4(new_n1345), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1341), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1339), .A2(new_n1344), .A3(new_n1354), .A4(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT61), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1357), .B1(new_n1340), .B2(new_n1326), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1359), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1360));
  AOI22_X1  g1160(.A1(new_n1266), .A2(G378), .B1(new_n1334), .B2(new_n1304), .ZN(new_n1361));
  NOR4_X1   g1161(.A1(new_n1361), .A2(KEYINPUT62), .A3(new_n1307), .A4(new_n1321), .ZN(new_n1362));
  NOR3_X1   g1162(.A1(new_n1358), .A2(new_n1360), .A3(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1356), .B1(new_n1363), .B2(new_n1354), .ZN(G405));
  AND2_X1   g1164(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1341), .A2(KEYINPUT127), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(G375), .A2(new_n1304), .ZN(new_n1368));
  AND2_X1   g1168(.A1(new_n1368), .A2(new_n1328), .ZN(new_n1369));
  AND2_X1   g1169(.A1(new_n1341), .A2(KEYINPUT127), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1370), .A2(new_n1354), .ZN(new_n1371));
  AND3_X1   g1171(.A1(new_n1367), .A2(new_n1369), .A3(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1369), .B1(new_n1367), .B2(new_n1371), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1372), .A2(new_n1373), .ZN(G402));
endmodule


