//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT91), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT16), .A3(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(G1gat), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT92), .B(G8gat), .Z(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT93), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(G8gat), .A3(new_n208), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215));
  XNOR2_X1  g014(.A(G57gat), .B(G64gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G71gat), .B(G78gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n214), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G231gat), .ZN(new_n224));
  INV_X1    g023(.A(G233gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n222), .B(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(G231gat), .A3(G233gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G211gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n215), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n240), .A3(new_n236), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(G29gat), .A2(G36gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT14), .ZN(new_n247));
  NAND2_X1  g046(.A1(G29gat), .A2(G36gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT89), .ZN(new_n249));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT15), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n250), .A2(KEYINPUT88), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n250), .B2(KEYINPUT88), .ZN(new_n253));
  AOI211_X1 g052(.A(new_n247), .B(new_n249), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n250), .ZN(new_n255));
  INV_X1    g054(.A(new_n247), .ZN(new_n256));
  AOI211_X1 g055(.A(new_n251), .B(new_n255), .C1(new_n256), .C2(new_n248), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  INV_X1    g059(.A(G85gat), .ZN(new_n261));
  INV_X1    g060(.A(G92gat), .ZN(new_n262));
  AOI22_X1  g061(.A1(KEYINPUT8), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT99), .ZN(new_n264));
  NAND2_X1  g063(.A1(G85gat), .A2(G92gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT7), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G99gat), .B(G106gat), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n267), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT90), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n258), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT17), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n245), .B(new_n271), .C1(new_n275), .C2(new_n270), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT100), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G190gat), .B(G218gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n279), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n269), .A3(new_n266), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT101), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(new_n220), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(new_n270), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n270), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G230gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(new_n225), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G120gat), .B(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(G176gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G204gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n270), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n288), .A2(new_n301), .A3(new_n289), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT102), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT102), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n304), .A3(new_n301), .A4(new_n289), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n300), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n293), .B(new_n299), .C1(new_n306), .C2(new_n292), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT103), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n306), .A2(new_n292), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n293), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n298), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n244), .A2(new_n283), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT98), .ZN(new_n315));
  AND2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  INV_X1    g116(.A(G169gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n295), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n227), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT65), .A4(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n324), .A2(new_n327), .A3(new_n326), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(new_n227), .A3(new_n325), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n324), .A3(new_n327), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n321), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n318), .A2(new_n295), .A3(KEYINPUT26), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(G169gat), .B2(G176gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n342), .B(new_n322), .C1(new_n344), .C2(new_n316), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n295), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT66), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n322), .A4(new_n342), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT27), .B(G183gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(new_n325), .ZN(new_n355));
  AND2_X1   g154(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n353), .B(new_n325), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n352), .A2(KEYINPUT67), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT67), .B1(new_n352), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n341), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G134gat), .ZN(new_n364));
  INV_X1    g163(.A(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G113gat), .ZN(new_n366));
  INV_X1    g165(.A(G113gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G120gat), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT1), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G127gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G113gat), .B(G120gat), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n372), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n364), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n370), .ZN(new_n375));
  OAI21_X1  g174(.A(G127gat), .B1(new_n372), .B2(KEYINPUT1), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(G134gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G227gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n225), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n375), .A2(new_n376), .A3(G134gat), .ZN(new_n383));
  AOI21_X1  g182(.A(G134gat), .B1(new_n375), .B2(new_n376), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n341), .C1(new_n361), .C2(new_n362), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT34), .ZN(new_n388));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n382), .B1(new_n379), .B2(new_n386), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(KEYINPUT33), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n386), .ZN(new_n397));
  AOI221_X4 g196(.A(new_n394), .B1(KEYINPUT33), .B2(new_n391), .C1(new_n397), .C2(new_n381), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n388), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT68), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n352), .A2(new_n360), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n352), .A2(new_n360), .A3(KEYINPUT67), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n385), .B1(new_n405), .B2(new_n341), .ZN(new_n406));
  INV_X1    g205(.A(new_n386), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n381), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n411), .A3(new_n391), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n395), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT34), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n387), .B(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT68), .B(new_n388), .C1(new_n396), .C2(new_n398), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT36), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n399), .A2(new_n416), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(KEYINPUT36), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n425), .A3(KEYINPUT36), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT70), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n329), .A2(new_n333), .B1(new_n339), .B2(new_n330), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n403), .B2(new_n404), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n432), .B2(KEYINPUT29), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT71), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT71), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n430), .C1(new_n432), .C2(KEYINPUT29), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n325), .B1(new_n356), .B2(new_n357), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT28), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n358), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n351), .B2(new_n346), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT72), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n341), .A2(new_n442), .A3(new_n401), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n443), .A3(new_n429), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n434), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(G197gat), .A2(G204gat), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT22), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G211gat), .A2(G218gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(G211gat), .A2(G218gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G218gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n232), .A2(new_n453), .A3(KEYINPUT22), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n449), .ZN(new_n455));
  XNOR2_X1  g254(.A(G197gat), .B(G204gat), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n448), .A2(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n445), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n430), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n448), .A2(new_n452), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT22), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n463), .A2(G211gat), .A3(G218gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n456), .B1(new_n464), .B2(new_n450), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n363), .A2(new_n429), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n461), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n458), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n471));
  XOR2_X1   g270(.A(G8gat), .B(G36gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G64gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(new_n262), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n468), .B1(new_n445), .B2(new_n457), .ZN(new_n476));
  INV_X1    g275(.A(new_n474), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT73), .B1(new_n476), .B2(new_n477), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  AND2_X1   g289(.A1(G155gat), .A2(G162gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(G155gat), .A2(G162gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G141gat), .B(G148gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT2), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(G155gat), .B2(G162gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G141gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G148gat), .ZN(new_n499));
  INV_X1    g298(.A(G148gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G141gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G155gat), .B(G162gat), .ZN(new_n503));
  INV_X1    g302(.A(G155gat), .ZN(new_n504));
  INV_X1    g303(.A(G162gat), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT2), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n385), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT79), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n507), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT3), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n378), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n509), .A2(KEYINPUT79), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(KEYINPUT79), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(KEYINPUT4), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G225gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT75), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n512), .A2(new_n517), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n511), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n385), .B2(new_n508), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n525), .B(new_n517), .C1(new_n526), .C2(new_n511), .ZN(new_n527));
  INV_X1    g326(.A(new_n522), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n378), .A2(new_n515), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n509), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n527), .B(KEYINPUT5), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(new_n483), .B(new_n490), .C1(new_n524), .C2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n490), .A3(new_n531), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n483), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n490), .B1(new_n524), .B2(new_n531), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n476), .A2(new_n477), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT74), .A4(new_n478), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n482), .A2(new_n537), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G78gat), .B(G106gat), .Z(new_n543));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n514), .A2(new_n459), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n457), .ZN(new_n546));
  INV_X1    g345(.A(G197gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n297), .ZN(new_n548));
  NAND2_X1  g347(.A1(G197gat), .A2(G204gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n463), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G211gat), .B(G218gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT81), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n448), .A2(new_n452), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n465), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT3), .B1(new_n555), .B2(new_n459), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n546), .B1(new_n556), .B2(new_n508), .ZN(new_n557));
  NAND2_X1  g356(.A1(G228gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT3), .B1(new_n466), .B2(new_n459), .ZN(new_n560));
  OAI211_X1 g359(.A(G228gat), .B(G233gat), .C1(new_n560), .C2(new_n508), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n466), .B1(new_n514), .B2(new_n459), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT82), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n513), .B1(new_n457), .B2(KEYINPUT29), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n564), .B2(new_n515), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT82), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n546), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G22gat), .ZN(new_n569));
  INV_X1    g368(.A(G22gat), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n559), .A2(new_n563), .A3(new_n570), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT80), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n544), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI211_X1 g373(.A(KEYINPUT80), .B(KEYINPUT31), .C1(new_n569), .C2(new_n571), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n543), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n466), .A2(new_n459), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n508), .B1(new_n577), .B2(new_n513), .ZN(new_n578));
  NOR4_X1   g377(.A1(new_n578), .A2(new_n562), .A3(KEYINPUT82), .A4(new_n558), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n566), .B1(new_n565), .B2(new_n546), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n570), .B1(new_n581), .B2(new_n559), .ZN(new_n582));
  AND4_X1   g381(.A1(new_n570), .A2(new_n559), .A3(new_n563), .A4(new_n567), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT31), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n572), .A2(new_n573), .A3(new_n544), .ZN(new_n586));
  INV_X1    g385(.A(new_n543), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT83), .B(G50gat), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n576), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n576), .B2(new_n588), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n542), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n427), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n512), .A2(new_n517), .A3(new_n520), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT85), .A3(new_n522), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT85), .B1(new_n597), .B2(new_n522), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n596), .B1(new_n526), .B2(new_n529), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n604), .A3(new_n490), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n540), .A2(new_n475), .A3(new_n478), .A4(new_n479), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n524), .A2(new_n531), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT86), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n524), .A2(KEYINPUT86), .A3(new_n531), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n490), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT40), .A4(new_n490), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n607), .A2(new_n608), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n534), .A2(new_n483), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n532), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n476), .B(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT38), .B1(new_n621), .B2(new_n477), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n445), .A2(new_n457), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n466), .B1(new_n461), .B2(new_n467), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n624), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n476), .A2(KEYINPUT37), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n623), .B(new_n474), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n619), .A2(new_n538), .A3(new_n622), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n592), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n617), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT84), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n427), .A2(new_n632), .A3(new_n593), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n595), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n490), .B1(new_n611), .B2(new_n612), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n533), .B1(new_n635), .B2(new_n535), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n636), .B(new_n423), .C1(new_n590), .C2(new_n591), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n637), .A2(KEYINPUT35), .A3(new_n608), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT87), .ZN(new_n640));
  INV_X1    g439(.A(new_n589), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n574), .A2(new_n575), .A3(new_n543), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n587), .B1(new_n585), .B2(new_n586), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n576), .A2(new_n588), .A3(new_n589), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n644), .A2(new_n645), .B1(new_n418), .B2(new_n417), .ZN(new_n646));
  INV_X1    g445(.A(new_n536), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n532), .B1(new_n618), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n481), .B2(new_n480), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n646), .A2(new_n540), .A3(new_n649), .A4(new_n541), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n640), .B1(new_n650), .B2(KEYINPUT35), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n419), .B1(new_n590), .B2(new_n591), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n640), .B(KEYINPUT35), .C1(new_n542), .C2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n639), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n634), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n273), .B(KEYINPUT17), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n214), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n212), .A2(new_n213), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT94), .B1(new_n275), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G229gat), .A2(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n259), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n659), .A2(new_n661), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT11), .B(G169gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G197gat), .ZN(new_n667));
  XOR2_X1   g466(.A(G113gat), .B(G141gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT12), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n212), .A2(new_n213), .A3(new_n258), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(KEYINPUT95), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n660), .A2(new_n674), .A3(new_n259), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n662), .B(KEYINPUT13), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n673), .A2(KEYINPUT96), .A3(new_n679), .A4(new_n675), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n670), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n664), .A2(KEYINPUT18), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n664), .A2(KEYINPUT18), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n685), .A2(new_n686), .B1(new_n678), .B2(new_n680), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n670), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n687), .A2(new_n683), .A3(new_n670), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n315), .B1(new_n656), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  AOI211_X1 g492(.A(KEYINPUT98), .B(new_n693), .C1(new_n634), .C2(new_n655), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n314), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n427), .A2(new_n632), .A3(new_n593), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n632), .B1(new_n427), .B2(new_n593), .ZN(new_n698));
  INV_X1    g497(.A(new_n631), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT35), .B1(new_n542), .B2(new_n652), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT87), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n638), .B1(new_n702), .B2(new_n653), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n691), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT98), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n656), .A2(new_n315), .A3(new_n691), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n314), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n696), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n648), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n608), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT16), .B(G8gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(G8gat), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(G1325gat));
  AOI21_X1  g518(.A(G15gat), .B1(new_n710), .B2(new_n423), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n427), .B1(new_n696), .B2(new_n709), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(G15gat), .B2(new_n721), .ZN(G1326gat));
  NAND2_X1  g521(.A1(new_n710), .A2(new_n592), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  INV_X1    g524(.A(new_n244), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n313), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n693), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n283), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n699), .A2(new_n594), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n702), .A2(new_n653), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n639), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT105), .B(new_n638), .C1(new_n702), .C2(new_n653), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT106), .B(new_n733), .C1(new_n736), .C2(new_n737), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n731), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n730), .B1(new_n656), .B2(new_n283), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n648), .B(new_n729), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G29gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n283), .B(new_n727), .C1(new_n692), .C2(new_n694), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n537), .ZN(new_n748));
  INV_X1    g547(.A(G29gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n747), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n537), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT107), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n745), .B(new_n754), .C1(new_n750), .C2(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1328gat));
  OAI211_X1 g555(.A(new_n608), .B(new_n729), .C1(new_n742), .C2(new_n743), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G36gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n728), .B1(new_n705), .B2(new_n706), .ZN(new_n759));
  INV_X1    g558(.A(G36gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n608), .A4(new_n283), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  INV_X1    g561(.A(new_n747), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n764), .A3(new_n760), .A4(new_n608), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n758), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT108), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n758), .A2(new_n765), .A3(new_n768), .A4(new_n762), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1329gat));
  INV_X1    g569(.A(new_n427), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(new_n729), .C1(new_n742), .C2(new_n743), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(G43gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n422), .A2(G43gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n763), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n774), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1330gat));
  NAND2_X1  g579(.A1(new_n747), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n707), .A2(new_n782), .A3(new_n283), .A4(new_n727), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n783), .A3(new_n592), .ZN(new_n784));
  INV_X1    g583(.A(G50gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n630), .A2(new_n785), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n729), .B(new_n787), .C1(new_n742), .C2(new_n743), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT48), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(new_n791), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1331gat));
  NAND2_X1  g592(.A1(new_n740), .A2(new_n741), .ZN(new_n794));
  INV_X1    g593(.A(new_n283), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n726), .A2(new_n693), .A3(new_n795), .A4(new_n313), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n648), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  INV_X1    g600(.A(new_n608), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  AND2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(G1333gat));
  NAND3_X1  g606(.A1(new_n799), .A2(G71gat), .A3(new_n771), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n798), .A2(new_n422), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(G71gat), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT50), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n808), .B(new_n812), .C1(G71gat), .C2(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1334gat));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n592), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT112), .B(G78gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1335gat));
  NOR2_X1   g616(.A1(new_n726), .A2(new_n691), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n738), .A2(new_n283), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n283), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(KEYINPUT113), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n822), .A2(new_n648), .A3(new_n313), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n742), .A2(new_n743), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n818), .A2(new_n313), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n648), .A2(G85gat), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n825), .A2(new_n261), .B1(new_n828), .B2(new_n830), .ZN(G1336gat));
  INV_X1    g630(.A(new_n827), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n608), .B(new_n832), .C1(new_n742), .C2(new_n743), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n833), .B2(G92gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n802), .A2(G92gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n822), .A2(new_n313), .A3(new_n824), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n312), .B1(new_n821), .B2(new_n823), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n833), .A2(G92gat), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(G1337gat));
  NAND2_X1  g640(.A1(new_n828), .A2(new_n771), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G99gat), .ZN(new_n843));
  INV_X1    g642(.A(G99gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n822), .A2(new_n844), .A3(new_n313), .A4(new_n824), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n422), .B2(new_n845), .ZN(G1338gat));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n822), .A2(new_n824), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n312), .A2(new_n630), .A3(G106gat), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT114), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n592), .B(new_n832), .C1(new_n742), .C2(new_n743), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(G106gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n850), .B1(new_n821), .B2(new_n823), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n852), .B2(G106gat), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n851), .A2(new_n853), .B1(new_n847), .B2(new_n855), .ZN(G1339gat));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n306), .B2(new_n292), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n309), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n306), .A2(new_n292), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n299), .B1(new_n860), .B2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n861), .A3(KEYINPUT55), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n308), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n689), .A2(new_n690), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n679), .B1(new_n673), .B2(new_n675), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT115), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(KEYINPUT115), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n869), .B(new_n870), .C1(new_n662), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n669), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n682), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n312), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n795), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(new_n866), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n283), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n726), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NOR4_X1   g678(.A1(new_n244), .A2(new_n691), .A3(new_n283), .A4(new_n313), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n608), .A2(new_n537), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n881), .A2(new_n652), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n367), .A3(new_n691), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n592), .A2(new_n422), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n886), .B(new_n882), .C1(new_n879), .C2(new_n880), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n691), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(G113gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n891), .B2(G113gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(G1340gat));
  NAND3_X1  g694(.A1(new_n884), .A2(new_n365), .A3(new_n313), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n889), .A2(new_n313), .A3(new_n890), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n365), .ZN(G1341gat));
  NAND4_X1  g697(.A1(new_n889), .A2(G127gat), .A3(new_n726), .A4(new_n890), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n884), .A2(new_n726), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(G127gat), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n901), .B(new_n902), .ZN(G1342gat));
  NOR2_X1   g702(.A1(new_n881), .A2(new_n883), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(new_n364), .A3(new_n646), .A4(new_n283), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT56), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n912), .A3(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n889), .A2(new_n283), .A3(new_n890), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT120), .B1(new_n915), .B2(G134gat), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n915), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n909), .B(new_n914), .C1(new_n916), .C2(new_n917), .ZN(G1343gat));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n919), .B(new_n592), .C1(new_n879), .C2(new_n880), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n771), .A2(new_n883), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT122), .Z(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n866), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT97), .B1(new_n687), .B2(new_n670), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n670), .B2(new_n687), .ZN(new_n926));
  INV_X1    g725(.A(new_n690), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n864), .A2(KEYINPUT123), .A3(new_n308), .A4(new_n865), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n924), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n875), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n283), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n878), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n244), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n314), .A2(new_n693), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n630), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n920), .B(new_n922), .C1(new_n935), .C2(new_n919), .ZN(new_n936));
  OAI21_X1  g735(.A(G141gat), .B1(new_n936), .B2(new_n693), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n881), .A2(new_n630), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n940), .A2(new_n498), .A3(new_n691), .A4(new_n921), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT58), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n937), .B(new_n941), .C1(new_n938), .C2(KEYINPUT58), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1344gat));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT57), .B1(new_n881), .B2(new_n630), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n935), .A2(new_n919), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n313), .A3(new_n922), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n951), .B2(G148gat), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n947), .B(G148gat), .C1(new_n936), .C2(new_n312), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n940), .A2(new_n921), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(new_n500), .A3(new_n313), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n958));
  OAI22_X1  g757(.A1(new_n952), .A2(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1345gat));
  AOI21_X1  g758(.A(G155gat), .B1(new_n955), .B2(new_n726), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n936), .A2(new_n504), .A3(new_n244), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1346gat));
  AOI21_X1  g761(.A(G162gat), .B1(new_n955), .B2(new_n283), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n936), .A2(new_n505), .A3(new_n795), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n881), .A2(new_n652), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n802), .A2(new_n648), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(new_n318), .A3(new_n691), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n967), .B(KEYINPUT126), .Z(new_n971));
  OAI211_X1 g770(.A(new_n886), .B(new_n971), .C1(new_n879), .C2(new_n880), .ZN(new_n972));
  OAI21_X1  g771(.A(G169gat), .B1(new_n972), .B2(new_n693), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n973), .ZN(G1348gat));
  NOR3_X1   g773(.A1(new_n972), .A2(new_n295), .A3(new_n312), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n969), .A2(new_n313), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n295), .ZN(G1349gat));
  OAI21_X1  g776(.A(G183gat), .B1(new_n972), .B2(new_n244), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n726), .A2(new_n354), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n968), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g780(.A1(new_n969), .A2(new_n325), .A3(new_n283), .ZN(new_n982));
  OAI21_X1  g781(.A(G190gat), .B1(new_n972), .B2(new_n795), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NAND3_X1  g785(.A1(new_n940), .A2(new_n427), .A3(new_n967), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(KEYINPUT127), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n988), .A2(new_n547), .A3(new_n691), .A4(new_n989), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n971), .A2(new_n427), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n950), .A2(new_n691), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n990), .B1(new_n547), .B2(new_n992), .ZN(G1352gat));
  NOR3_X1   g792(.A1(new_n987), .A2(G204gat), .A3(new_n312), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n950), .A2(new_n313), .A3(new_n991), .ZN(new_n998));
  OAI211_X1 g797(.A(new_n996), .B(new_n997), .C1(new_n297), .C2(new_n998), .ZN(G1353gat));
  NAND4_X1  g798(.A1(new_n988), .A2(new_n232), .A3(new_n726), .A4(new_n989), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n950), .A2(new_n726), .A3(new_n991), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(G211gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G1354gat));
  NAND4_X1  g803(.A1(new_n988), .A2(new_n453), .A3(new_n283), .A4(new_n989), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n950), .A2(new_n283), .A3(new_n991), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n453), .B2(new_n1006), .ZN(G1355gat));
endmodule


