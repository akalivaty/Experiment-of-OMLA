//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT2), .A2(G113), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT68), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT2), .A2(G113), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(G116), .B(G119), .Z(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G116), .B(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n190), .A2(new_n197), .A3(new_n193), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G104), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n205), .A2(G107), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(new_n203), .ZN(new_n211));
  INV_X1    g025(.A(new_n201), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n207), .A4(new_n206), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n209), .A3(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(new_n210), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n201), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G116), .ZN(new_n223));
  OAI211_X1 g037(.A(G113), .B(new_n223), .C1(new_n195), .C2(new_n221), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n198), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n217), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT6), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n227), .B1(new_n217), .B2(new_n226), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI211_X1 g045(.A(KEYINPUT6), .B(new_n227), .C1(new_n217), .C2(new_n226), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT64), .A2(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(G143), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(G143), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT64), .A2(G146), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT64), .A2(G146), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n247), .B2(G143), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n242), .A2(new_n243), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G125), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n241), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n258));
  INV_X1    g072(.A(new_n244), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT64), .B(G146), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(new_n239), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n256), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n253), .B1(new_n247), .B2(G143), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT67), .B(new_n248), .C1(new_n263), .C2(new_n257), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n255), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n252), .B1(new_n265), .B2(G125), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G224), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT84), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(G902), .B1(new_n233), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n227), .B(KEYINPUT8), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n220), .A2(new_n225), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n226), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n266), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(KEYINPUT7), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT86), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT7), .B1(new_n268), .B2(KEYINPUT85), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(KEYINPUT85), .B2(new_n268), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n266), .B2(new_n280), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n277), .B(KEYINPUT87), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n228), .ZN(new_n285));
  INV_X1    g099(.A(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT87), .B1(new_n287), .B2(new_n277), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n271), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n277), .B1(new_n282), .B2(new_n283), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n284), .A3(new_n228), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n290), .A3(new_n271), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n188), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT9), .B(G234), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT80), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT94), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n306));
  XNOR2_X1  g120(.A(G113), .B(G122), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT92), .B(G104), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(KEYINPUT88), .A2(G143), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT88), .A2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G237), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n313), .A2(new_n267), .A3(G214), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G131), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n267), .A3(G214), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n311), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT91), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n315), .A2(new_n318), .A3(new_n321), .A4(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n331), .A3(KEYINPUT76), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n326), .A2(KEYINPUT76), .A3(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n329), .B1(new_n334), .B2(new_n328), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G146), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(KEYINPUT90), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(KEYINPUT19), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n327), .A2(new_n331), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(KEYINPUT19), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n325), .B(new_n336), .C1(new_n342), .C2(new_n260), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n317), .B1(new_n310), .B2(new_n311), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n317), .A2(new_n311), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT18), .A2(G131), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT89), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT89), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n323), .A2(new_n349), .A3(KEYINPUT18), .A4(G131), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n337), .A2(G146), .A3(new_n339), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n327), .A2(new_n331), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n247), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n346), .A2(new_n347), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n309), .B1(new_n343), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n320), .A2(new_n324), .A3(new_n359), .A4(new_n322), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n335), .A2(G146), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n323), .A2(KEYINPUT17), .A3(G131), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n336), .A4(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n357), .A3(new_n309), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT93), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n363), .A2(new_n357), .A3(KEYINPUT93), .A4(new_n309), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n358), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G475), .ZN(new_n369));
  INV_X1    g183(.A(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n305), .B(new_n306), .C1(new_n368), .C2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n309), .B1(new_n363), .B2(new_n357), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n366), .B2(new_n367), .ZN(new_n374));
  OAI21_X1  g188(.A(G475), .B1(new_n374), .B2(G902), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n366), .A2(new_n367), .ZN(new_n377));
  INV_X1    g191(.A(new_n358), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n379), .A2(KEYINPUT94), .A3(new_n369), .A4(new_n370), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n305), .B1(new_n368), .B2(new_n371), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(KEYINPUT20), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n267), .A2(G952), .ZN(new_n383));
  INV_X1    g197(.A(G234), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n313), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT21), .B(G898), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT97), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n370), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G478), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G116), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT14), .A3(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(G116), .B(G122), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(G107), .B(new_n396), .C1(new_n398), .C2(KEYINPUT14), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n200), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT65), .B(G134), .ZN(new_n401));
  XNOR2_X1  g215(.A(G128), .B(G143), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n401), .A2(new_n402), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n399), .B(new_n400), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(KEYINPUT13), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n239), .A2(G128), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n407), .B(G134), .C1(KEYINPUT13), .C2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n397), .B(new_n200), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n403), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n267), .A2(G217), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n301), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n411), .A3(new_n414), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n406), .A2(new_n414), .A3(new_n411), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n406), .B2(new_n411), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n419), .B(new_n370), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n394), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n393), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n370), .B1(new_n421), .B2(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT95), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n393), .B1(new_n430), .B2(new_n423), .ZN(new_n431));
  INV_X1    g245(.A(new_n427), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT96), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n391), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n376), .A2(new_n382), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G469), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT12), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n265), .A2(new_n438), .A3(new_n220), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT11), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n401), .B2(G137), .ZN(new_n441));
  INV_X1    g255(.A(G134), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G137), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n401), .B2(G137), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G131), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n316), .B(new_n441), .C1(new_n444), .C2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n257), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n238), .B2(new_n240), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n215), .B(new_n219), .C1(new_n255), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n265), .B2(new_n220), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n437), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n265), .A2(new_n220), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT83), .A3(new_n452), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n457), .A2(KEYINPUT12), .A3(new_n448), .A4(new_n439), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n210), .A2(new_n251), .A3(new_n216), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n452), .A2(KEYINPUT82), .A3(new_n461), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n255), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n245), .A2(new_n246), .A3(new_n239), .ZN(new_n468));
  OAI21_X1  g282(.A(G128), .B1(new_n468), .B2(new_n253), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT67), .B1(new_n469), .B2(new_n248), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n258), .A2(new_n261), .A3(new_n256), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n265), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n220), .A2(new_n461), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n466), .A2(new_n446), .A3(new_n477), .A4(new_n447), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G140), .ZN(new_n479));
  INV_X1    g293(.A(G227), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n479), .B(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n459), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n477), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n448), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n487), .B2(new_n478), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n436), .B(new_n370), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n478), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n482), .B1(new_n459), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n478), .A3(new_n483), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(G469), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n436), .A2(new_n370), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AND4_X1   g310(.A1(new_n298), .A2(new_n304), .A3(new_n435), .A4(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G217), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(G234), .B2(new_n370), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G137), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n361), .A2(new_n336), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n222), .A2(G128), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT75), .B1(new_n257), .B2(G119), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n507), .B(new_n508), .Z(new_n509));
  INV_X1    g323(.A(G110), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n257), .A2(G119), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT24), .B(G110), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n505), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT77), .B(G110), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n354), .B(new_n336), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n504), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n519), .A3(new_n504), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n501), .B1(new_n523), .B2(G902), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n521), .A2(KEYINPUT25), .A3(new_n370), .A4(new_n522), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n500), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n523), .A2(G902), .A3(new_n499), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n313), .A2(new_n267), .A3(G210), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT27), .Z(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT26), .B(G101), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n531), .B(new_n532), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n401), .A2(G137), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n442), .A2(G137), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n447), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n473), .A2(new_n475), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n448), .A2(new_n251), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT71), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n199), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT72), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n539), .A2(new_n545), .A3(new_n540), .A4(new_n542), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n447), .A2(KEYINPUT66), .A3(new_n537), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT66), .B1(new_n447), .B2(new_n537), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n547), .A2(new_n265), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n540), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n199), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n544), .A2(new_n546), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n539), .A2(KEYINPUT30), .A3(new_n540), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n549), .B2(new_n550), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n199), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n557), .A2(KEYINPUT31), .A3(new_n561), .A4(new_n533), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n544), .A3(new_n546), .A4(new_n533), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n534), .A2(new_n556), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT73), .B1(G472), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(KEYINPUT73), .A2(G472), .A3(G902), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT32), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n563), .A2(new_n564), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n563), .A2(new_n564), .ZN(new_n573));
  INV_X1    g387(.A(new_n555), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n552), .B2(KEYINPUT28), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n572), .A2(new_n573), .B1(new_n533), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT32), .ZN(new_n577));
  INV_X1    g391(.A(new_n570), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n557), .A2(new_n561), .A3(new_n534), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n575), .B2(new_n534), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT29), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n539), .A2(new_n540), .ZN(new_n585));
  INV_X1    g399(.A(new_n542), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n589), .A3(new_n586), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n588), .A2(new_n544), .A3(new_n546), .A4(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n574), .B1(new_n591), .B2(KEYINPUT28), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n534), .A2(new_n583), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n529), .B1(new_n580), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT78), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n571), .A2(new_n579), .B1(new_n595), .B2(G472), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(KEYINPUT78), .A3(new_n529), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n497), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT98), .B(G101), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n576), .B2(new_n370), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n566), .A2(new_n570), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n496), .A2(new_n304), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n529), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n376), .A2(new_n382), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n416), .A2(new_n417), .B1(new_n613), .B2(KEYINPUT33), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(KEYINPUT33), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n614), .B(new_n615), .Z(new_n616));
  NOR2_X1   g430(.A1(new_n392), .A2(G902), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n616), .A2(new_n617), .B1(new_n392), .B2(new_n429), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n391), .ZN(new_n621));
  INV_X1    g435(.A(new_n297), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n290), .B1(new_n296), .B2(new_n271), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n187), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n611), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT100), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND2_X1  g442(.A1(new_n372), .A2(new_n375), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n368), .A2(new_n371), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n306), .B1(new_n630), .B2(KEYINPUT94), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n631), .B2(new_n381), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n428), .A2(new_n433), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n624), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n608), .A2(new_n635), .A3(new_n610), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NAND2_X1  g452(.A1(new_n515), .A2(new_n519), .ZN(new_n639));
  INV_X1    g453(.A(new_n504), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n639), .B1(KEYINPUT36), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n499), .A2(G902), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(KEYINPUT36), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n515), .A2(new_n519), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n526), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n497), .A2(new_n608), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  NAND3_X1  g464(.A1(new_n298), .A2(new_n304), .A3(new_n496), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n647), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n386), .B1(new_n390), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n376), .A2(new_n382), .A3(new_n633), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n556), .A2(new_n534), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n562), .A2(new_n565), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT32), .B(new_n570), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n605), .B1(new_n584), .B2(new_n594), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n652), .B(new_n658), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  NAND2_X1  g480(.A1(new_n557), .A2(new_n561), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n533), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n370), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n591), .A2(new_n533), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n661), .B2(new_n662), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n622), .A2(new_n623), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT102), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n673), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n428), .A2(new_n433), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n376), .B2(new_n382), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n647), .A2(new_n188), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n672), .A2(new_n676), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n609), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n655), .B(KEYINPUT39), .Z(new_n682));
  AOI21_X1  g496(.A(KEYINPUT104), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n681), .A2(KEYINPUT104), .A3(new_n682), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n686), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT40), .B1(new_n688), .B2(new_n683), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n680), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n680), .A2(new_n692), .A3(new_n689), .A4(new_n687), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n239), .ZN(G45));
  AOI21_X1  g509(.A(new_n618), .B1(new_n376), .B2(new_n382), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n656), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n653), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n652), .B(new_n698), .C1(new_n663), .C2(new_n664), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NAND2_X1  g514(.A1(new_n580), .A2(new_n596), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n624), .A2(new_n620), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n485), .A2(new_n488), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n436), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n370), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n370), .B1(new_n485), .B2(new_n488), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n705), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n304), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n701), .A2(new_n528), .A3(new_n702), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n701), .A2(new_n528), .A3(new_n635), .A4(new_n711), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NAND2_X1  g530(.A1(new_n647), .A2(new_n435), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n292), .A2(new_n297), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n187), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n717), .A2(new_n719), .A3(new_n710), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n701), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  XOR2_X1   g536(.A(new_n570), .B(KEYINPUT107), .Z(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n589), .B1(new_n585), .B2(new_n586), .ZN(new_n725));
  AOI211_X1 g539(.A(KEYINPUT74), .B(new_n542), .C1(new_n539), .C2(new_n540), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n554), .B1(new_n557), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n534), .B1(new_n728), .B2(new_n574), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n724), .B1(new_n729), .B2(new_n660), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n606), .A2(new_n730), .A3(new_n529), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n298), .A2(new_n678), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n707), .A2(new_n709), .A3(new_n304), .A4(new_n621), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR3_X1   g550(.A1(new_n719), .A2(new_n697), .A3(new_n710), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n606), .A2(new_n653), .A3(new_n730), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  INV_X1    g554(.A(new_n697), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n493), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n491), .A2(KEYINPUT108), .A3(G469), .A4(new_n492), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n489), .A3(new_n495), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n673), .A3(new_n187), .A4(new_n304), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n701), .A2(new_n528), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n597), .A2(KEYINPUT42), .A3(new_n741), .A4(new_n747), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n316), .ZN(G33));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n632), .A2(new_n756), .A3(new_n633), .A4(new_n656), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n657), .A2(KEYINPUT109), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n600), .A2(new_n529), .A3(new_n746), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n442), .ZN(G36));
  AOI21_X1  g575(.A(KEYINPUT113), .B1(new_n632), .B2(new_n619), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT43), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n632), .A2(new_n619), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n608), .A3(new_n653), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n718), .A2(new_n188), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n491), .A2(new_n492), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n436), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT110), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n774), .B2(KEYINPUT110), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n494), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT111), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n489), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n304), .A3(new_n682), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(KEYINPUT112), .A3(new_n304), .A4(new_n682), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n771), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  AND4_X1   g605(.A1(new_n600), .A2(new_n529), .A3(new_n741), .A4(new_n770), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n304), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT47), .B1(new_n784), .B2(new_n304), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  INV_X1    g610(.A(new_n767), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n386), .A3(new_n711), .A4(new_n770), .ZN(new_n798));
  INV_X1    g612(.A(new_n730), .ZN(new_n799));
  OAI21_X1  g613(.A(G472), .B1(new_n566), .B2(G902), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n798), .A2(new_n653), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n672), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n529), .A2(new_n385), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n711), .A3(new_n770), .A4(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n612), .A3(new_n619), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n676), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n711), .A3(new_n188), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT120), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n797), .A2(new_n386), .A3(new_n731), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n809), .B(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n812), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT50), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n707), .A2(new_n709), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n304), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n793), .A2(new_n794), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n770), .ZN(new_n821));
  OAI221_X1 g635(.A(new_n807), .B1(new_n813), .B2(new_n817), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n597), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n798), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n812), .A2(new_n719), .A3(new_n710), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n383), .B1(new_n805), .B2(new_n620), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n824), .B(new_n830), .C1(new_n832), .C2(new_n823), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n425), .A2(new_n427), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n655), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n632), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n632), .A2(KEYINPUT117), .A3(new_n835), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n681), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n741), .A2(new_n304), .A3(new_n745), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n600), .A2(new_n840), .B1(new_n841), .B2(new_n801), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n653), .A2(new_n188), .A3(new_n718), .ZN(new_n843));
  AOI221_X4 g657(.A(new_n760), .B1(new_n842), .B2(new_n843), .C1(new_n750), .C2(new_n752), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n701), .A2(new_n720), .B1(new_n731), .B2(new_n734), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n712), .A3(new_n715), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n712), .A3(new_n715), .A4(KEYINPUT114), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT115), .B1(new_n624), .B2(new_n620), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n298), .A2(new_n852), .A3(new_n696), .A4(new_n621), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(new_n608), .A3(new_n610), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n376), .A2(new_n382), .A3(new_n834), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n624), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n608), .A2(new_n857), .A3(new_n858), .A4(new_n610), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(new_n859), .A3(new_n648), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT78), .B1(new_n600), .B2(new_n529), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n701), .A2(new_n598), .A3(new_n528), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n863), .B2(new_n497), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n844), .A2(new_n850), .A3(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n526), .A2(new_n646), .A3(new_n655), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n298), .A2(new_n866), .A3(new_n678), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n745), .A2(new_n304), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n672), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n665), .A2(new_n699), .A3(new_n739), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n651), .B1(new_n580), .B2(new_n596), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n874), .A2(new_n658), .B1(new_n738), .B2(new_n737), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n699), .A4(new_n870), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n865), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n860), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n602), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n848), .B2(new_n849), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n873), .A2(new_n876), .A3(KEYINPUT118), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n884), .A3(new_n844), .A4(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n879), .A2(KEYINPUT53), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n885), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n890), .B2(new_n865), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  INV_X1    g706(.A(new_n846), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n864), .A2(new_n893), .A3(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n842), .A2(new_n843), .ZN(new_n895));
  INV_X1    g709(.A(new_n760), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n895), .B(new_n896), .C1(new_n751), .C2(new_n753), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n878), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n892), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n889), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n833), .A2(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n818), .A2(KEYINPUT49), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n818), .A2(KEYINPUT49), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n528), .A2(new_n187), .A3(new_n304), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n764), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n803), .A3(new_n808), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n907), .ZN(G75));
  AOI21_X1  g722(.A(new_n898), .B1(new_n886), .B2(new_n887), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n370), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n233), .B(new_n270), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n911), .B2(new_n912), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n267), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  INV_X1    g732(.A(new_n887), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n844), .A2(new_n850), .A3(new_n864), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n873), .A2(new_n876), .A3(KEYINPUT118), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT118), .B1(new_n873), .B2(new_n876), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT54), .B1(new_n924), .B2(new_n898), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n900), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT122), .B(KEYINPUT54), .C1(new_n924), .C2(new_n898), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n494), .B(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n703), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n910), .A2(new_n775), .A3(new_n777), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n917), .B1(new_n931), .B2(new_n932), .ZN(G54));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n910), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT123), .B1(new_n935), .B2(new_n368), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n917), .B1(new_n935), .B2(new_n368), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n910), .A2(new_n938), .A3(new_n379), .A4(new_n934), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(G60));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT59), .Z(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n889), .B2(new_n900), .ZN(new_n943));
  OAI22_X1  g757(.A1(new_n943), .A2(new_n616), .B1(G952), .B2(new_n267), .ZN(new_n944));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n616), .A2(new_n927), .A3(new_n928), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n924), .B2(new_n898), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n917), .B1(new_n951), .B2(new_n523), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n891), .B2(new_n899), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n641), .A2(new_n644), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR4_X1   g771(.A1(new_n909), .A2(KEYINPUT124), .A3(new_n955), .A4(new_n949), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n952), .B(KEYINPUT61), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  AOI21_X1  g777(.A(new_n267), .B1(new_n388), .B2(G224), .ZN(new_n964));
  INV_X1    g778(.A(new_n882), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n267), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT125), .ZN(new_n967));
  OAI22_X1  g781(.A1(new_n231), .A2(new_n232), .B1(G898), .B2(new_n267), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  NAND2_X1  g783(.A1(new_n558), .A2(new_n560), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT126), .Z(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(new_n342), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n875), .A2(new_n699), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n691), .A2(new_n693), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n688), .A2(new_n683), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n857), .A2(new_n696), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n863), .A2(new_n978), .A3(new_n770), .A4(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n977), .A2(new_n790), .A3(new_n795), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n973), .B1(new_n981), .B2(new_n267), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n480), .B2(new_n654), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT127), .B1(new_n790), .B2(new_n974), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n790), .A2(KEYINPUT127), .A3(new_n974), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n825), .A2(new_n732), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n787), .A2(new_n788), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n754), .A2(new_n760), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n990), .A2(new_n795), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n973), .A2(new_n267), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n983), .B(new_n984), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n988), .B2(new_n992), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n996), .A2(new_n982), .A3(new_n654), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n997), .B2(new_n984), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n981), .B2(new_n965), .ZN(new_n1001));
  INV_X1    g815(.A(new_n668), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n668), .A2(new_n581), .A3(new_n1000), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n917), .B1(new_n888), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n581), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n988), .A2(new_n992), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1000), .B1(new_n1008), .B2(new_n965), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(G57));
endmodule


