//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  AND4_X1   g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT66), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT67), .Z(new_n218));
  INV_X1    g0018(.A(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(new_n215), .A2(new_n216), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g0032(.A1(new_n218), .A2(new_n223), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n228), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n224), .ZN(new_n253));
  INV_X1    g0053(.A(G107), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n254), .A2(KEYINPUT23), .A3(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT23), .B1(new_n254), .B2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G116), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n255), .A2(new_n256), .B1(G20), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n225), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT22), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT22), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n263), .A2(new_n264), .A3(new_n225), .A4(G87), .ZN(new_n265));
  AOI211_X1 g0065(.A(KEYINPUT24), .B(new_n258), .C1(new_n262), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT24), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(new_n258), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(KEYINPUT84), .B(new_n253), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n253), .B1(new_n266), .B2(new_n270), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT84), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n225), .A2(G107), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n219), .A2(G1), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT85), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT25), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n278), .A2(KEYINPUT25), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(KEYINPUT25), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(new_n275), .A3(new_n276), .A4(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n252), .A2(new_n224), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n276), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n283), .B(new_n284), .C1(G1), .C2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n279), .B(new_n282), .C1(new_n286), .C2(new_n254), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  OAI211_X1 g0090(.A(G250), .B(new_n290), .C1(new_n259), .C2(new_n260), .ZN(new_n291));
  INV_X1    g0091(.A(G294), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n289), .B(new_n291), .C1(new_n285), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G1), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT5), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT5), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G264), .ZN(new_n306));
  INV_X1    g0106(.A(G1), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(G45), .C1(new_n298), .C2(KEYINPUT5), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT79), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G274), .ZN(new_n311));
  INV_X1    g0111(.A(new_n224), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n303), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n297), .A2(KEYINPUT79), .A3(new_n301), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n313), .A3(new_n314), .A4(new_n299), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n295), .A2(new_n306), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n293), .A2(new_n294), .B1(new_n305), .B2(G264), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  AND4_X1   g0122(.A1(new_n271), .A2(new_n274), .A3(new_n288), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G179), .B2(new_n316), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n287), .B1(new_n272), .B2(new_n273), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n271), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n219), .A2(new_n225), .A3(G1), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n228), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT12), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G20), .A2(G33), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(G50), .B1(G20), .B2(new_n228), .ZN(new_n334));
  INV_X1    g0134(.A(G77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n225), .A2(G33), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n283), .A2(new_n284), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n307), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G68), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n332), .B(new_n338), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT11), .B1(new_n337), .B2(new_n253), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  INV_X1    g0146(.A(G226), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n290), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n235), .A2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(new_n349), .C1(new_n259), .C2(new_n260), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n304), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g0154(.A(KEYINPUT71), .B(new_n304), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n307), .B1(G41), .B2(G45), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(new_n304), .A3(G274), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n304), .A2(G238), .A3(new_n356), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT72), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT72), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n354), .A2(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G226), .A2(G1698), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n235), .B2(G1698), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n263), .B1(G33), .B2(G97), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT71), .B1(new_n367), .B2(new_n304), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n352), .A2(new_n353), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n358), .A2(new_n359), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n364), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n346), .B(G169), .C1(new_n363), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n375), .A3(new_n364), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(G179), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n346), .B1(new_n382), .B2(G169), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n345), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G200), .B1(new_n363), .B2(new_n376), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(G190), .A3(new_n379), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n344), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n388), .B(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n204), .A2(G20), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT8), .B(G58), .ZN(new_n392));
  INV_X1    g0192(.A(G150), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n225), .A2(new_n285), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n392), .A2(new_n336), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n253), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n340), .A2(G50), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n339), .A2(new_n397), .B1(G50), .B2(new_n284), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(new_n400), .B(KEYINPUT9), .Z(new_n401));
  OR2_X1    g0201(.A1(KEYINPUT3), .A2(G33), .ZN(new_n402));
  NAND2_X1  g0202(.A1(KEYINPUT3), .A2(G33), .ZN(new_n403));
  AOI21_X1  g0203(.A(G1698), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G222), .ZN(new_n405));
  INV_X1    g0205(.A(G223), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n263), .A2(G1698), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n405), .B1(new_n335), .B2(new_n263), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n294), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n304), .A2(new_n356), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(G226), .B1(new_n313), .B2(new_n357), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G200), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n320), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT10), .B1(new_n401), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n400), .B(KEYINPUT9), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n414), .A2(KEYINPUT70), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n409), .A2(new_n412), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT10), .B1(new_n419), .B2(G190), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(KEYINPUT70), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n417), .A2(new_n418), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n400), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n413), .B2(new_n324), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT68), .B(G179), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  INV_X1    g0227(.A(G244), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n358), .B1(new_n428), .B2(new_n410), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT69), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  INV_X1    g0232(.A(G238), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n407), .A2(new_n433), .B1(new_n254), .B2(new_n263), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(G232), .B2(new_n404), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n431), .B(new_n432), .C1(new_n435), .C2(new_n304), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n436), .A2(new_n426), .ZN(new_n437));
  INV_X1    g0237(.A(new_n392), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n333), .B1(G20), .B2(G77), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(new_n336), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n283), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n340), .A2(G77), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n339), .A2(new_n443), .B1(G77), .B2(new_n284), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n436), .A2(new_n324), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n437), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n436), .B2(G200), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n320), .B2(new_n436), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n423), .A2(new_n427), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n438), .A2(new_n340), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n452), .A2(new_n339), .B1(new_n284), .B2(new_n438), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n347), .A2(G1698), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n263), .B(new_n455), .C1(G223), .C2(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n294), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n358), .B1(new_n235), .B2(new_n410), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(G200), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n304), .B1(new_n456), .B2(new_n457), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n463), .A2(new_n460), .A3(G190), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT75), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n402), .A2(new_n225), .A3(new_n403), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT7), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n259), .A2(new_n260), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G68), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G58), .A2(G68), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n225), .B1(new_n229), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G159), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n394), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT74), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(G58), .A2(G68), .ZN(new_n480));
  OAI21_X1  g0280(.A(G20), .B1(new_n480), .B2(new_n201), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT74), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n333), .A2(G159), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT16), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n283), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n474), .A2(KEYINPUT16), .A3(new_n485), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n467), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n228), .B1(new_n470), .B2(new_n472), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(new_n489), .A3(new_n467), .A4(new_n253), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n454), .B(new_n466), .C1(new_n490), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT17), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n498), .B(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n454), .B1(new_n490), .B2(new_n497), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT18), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n463), .A2(new_n460), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n426), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n324), .B2(new_n503), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n473), .A2(G68), .B1(new_n479), .B2(new_n484), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n253), .B1(new_n507), .B2(KEYINPUT16), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n493), .A2(new_n494), .A3(new_n487), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT75), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n453), .B1(new_n510), .B2(new_n496), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n503), .A2(new_n324), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n426), .B2(new_n503), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT18), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n500), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n390), .A2(new_n451), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n286), .A2(G116), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G116), .B2(new_n330), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n225), .C1(G33), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT20), .ZN(new_n524));
  INV_X1    g0324(.A(G116), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(G20), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n526), .A3(new_n253), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n300), .A2(G41), .ZN(new_n531));
  OAI211_X1 g0331(.A(G270), .B(new_n304), .C1(new_n308), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT82), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT82), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n302), .A2(new_n534), .A3(G270), .A4(new_n304), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n537));
  OAI211_X1 g0337(.A(G257), .B(new_n290), .C1(new_n259), .C2(new_n260), .ZN(new_n538));
  INV_X1    g0338(.A(G303), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n263), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n294), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(new_n541), .A3(new_n315), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(new_n320), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n530), .B(new_n543), .C1(G200), .C2(new_n542), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n530), .A2(G169), .A3(new_n542), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n536), .A2(new_n541), .A3(G179), .A4(new_n315), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n530), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n530), .A2(KEYINPUT21), .A3(G169), .A4(new_n542), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n225), .B1(new_n351), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G87), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n521), .A3(new_n254), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n225), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n336), .B2(new_n521), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n253), .B1(new_n330), .B2(new_n440), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n286), .B2(new_n440), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n433), .A2(new_n290), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n428), .A2(G1698), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n259), .C2(new_n260), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n304), .B1(new_n566), .B2(new_n257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n297), .A2(new_n311), .ZN(new_n568));
  INV_X1    g0368(.A(G250), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n296), .B2(G1), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n568), .A2(new_n304), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(G169), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n304), .A3(new_n570), .ZN(new_n573));
  INV_X1    g0373(.A(new_n257), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G238), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n428), .B2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(new_n263), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n426), .B(new_n573), .C1(new_n577), .C2(new_n304), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n563), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n567), .B2(new_n571), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n286), .A2(new_n556), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n562), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G190), .B(new_n573), .C1(new_n577), .C2(new_n304), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n567), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(KEYINPUT80), .A3(G190), .A4(new_n573), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT81), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n580), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(new_n290), .C1(new_n259), .C2(new_n260), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n428), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n263), .A2(new_n290), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n520), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G250), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n263), .A2(KEYINPUT78), .A3(G250), .A4(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n294), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n426), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n302), .A2(G257), .A3(new_n304), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n315), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n324), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n254), .B1(new_n470), .B2(new_n472), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n394), .A2(new_n335), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n521), .A2(new_n254), .A3(KEYINPUT6), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G97), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n254), .A2(KEYINPUT76), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT76), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G107), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n615), .A2(new_n617), .A3(new_n619), .A4(new_n621), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n614), .B1(new_n625), .B2(G20), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n613), .B1(new_n626), .B2(KEYINPUT77), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT77), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n225), .B1(new_n623), .B2(new_n624), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n614), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n283), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n330), .A2(new_n521), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n286), .B2(new_n521), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n610), .B(new_n612), .C1(new_n631), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n625), .A2(G20), .ZN(new_n635));
  INV_X1    g0435(.A(new_n614), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(KEYINPUT77), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n613), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n630), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n639), .B2(new_n253), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n605), .A2(new_n320), .A3(new_n609), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n404), .A2(new_n597), .B1(G33), .B2(G283), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n596), .A3(new_n602), .A4(new_n603), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n608), .B1(new_n643), .B2(new_n294), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n644), .B2(G200), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n593), .A2(new_n634), .A3(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n329), .A2(new_n517), .A3(new_n553), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n427), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n502), .B1(new_n501), .B2(new_n505), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n511), .A2(KEYINPUT18), .A3(new_n513), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n506), .A2(new_n514), .A3(KEYINPUT89), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n448), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n387), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n657), .A2(new_n384), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n500), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n423), .A2(KEYINPUT90), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT90), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n416), .A2(new_n422), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n649), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n517), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n612), .A2(new_n610), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n640), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n666), .A2(new_n668), .A3(new_n593), .A4(KEYINPUT26), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT87), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n583), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n562), .A2(new_n581), .A3(new_n582), .A4(KEYINPUT87), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n589), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n572), .A2(new_n578), .A3(KEYINPUT86), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT86), .B1(new_n572), .B2(new_n578), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n563), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n634), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n666), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n668), .A2(new_n593), .A3(KEYINPUT26), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n327), .A2(new_n271), .A3(new_n322), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n634), .A3(new_n646), .A4(new_n673), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n328), .A2(new_n552), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n664), .B1(new_n665), .B2(new_n686), .ZN(G369));
  INV_X1    g0487(.A(new_n530), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n276), .A2(new_n225), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n553), .B1(new_n688), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n552), .A2(new_n530), .A3(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n328), .A2(new_n694), .ZN(new_n702));
  INV_X1    g0502(.A(new_n329), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n695), .B1(new_n327), .B2(new_n271), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT91), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n552), .A2(new_n695), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(new_n329), .B1(new_n328), .B2(new_n695), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(G399));
  NOR2_X1   g0511(.A1(new_n220), .A2(G41), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n557), .A2(G116), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n712), .A2(new_n307), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n231), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NOR3_X1   g0516(.A1(new_n686), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT26), .B1(new_n634), .B2(new_n677), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n668), .A2(new_n593), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT26), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n695), .B1(new_n685), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n647), .A2(new_n329), .A3(new_n553), .A4(new_n695), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT92), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n567), .A2(new_n571), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n605), .A2(new_n319), .A3(new_n609), .A4(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n729), .B2(new_n548), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n728), .A2(new_n295), .A3(new_n306), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n549), .A2(new_n644), .A3(KEYINPUT30), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n728), .A2(new_n426), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n611), .A2(new_n316), .A3(new_n542), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n735), .B2(new_n694), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n726), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(new_n726), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n725), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n724), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n716), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(new_n712), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n219), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n307), .B1(new_n746), .B2(G45), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(KEYINPUT93), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT93), .ZN(new_n749));
  INV_X1    g0549(.A(new_n747), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n749), .B1(new_n712), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n699), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n224), .B1(G20), .B2(new_n324), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n225), .A2(G190), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT95), .B(G159), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT32), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n225), .A2(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n225), .A2(new_n317), .A3(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n426), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G68), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n426), .A2(new_n758), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n765), .A2(new_n320), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n777), .A2(G77), .B1(new_n779), .B2(G107), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n764), .A2(new_n771), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n320), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n225), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n471), .B1(new_n784), .B2(G97), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n225), .A2(new_n320), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n426), .A2(G200), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n426), .A2(new_n317), .A3(new_n786), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n785), .B1(new_n787), .B2(new_n202), .C1(new_n227), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n263), .B1(new_n784), .B2(G294), .ZN(new_n790));
  INV_X1    g0590(.A(G326), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(new_n787), .B2(new_n791), .C1(new_n792), .C2(new_n788), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n774), .A2(new_n794), .B1(G283), .B2(new_n779), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n777), .A2(G311), .B1(new_n761), .B2(G329), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(new_n769), .C2(new_n539), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n781), .A2(new_n789), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n220), .A2(new_n471), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n525), .B2(new_n220), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n221), .A2(new_n471), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n231), .A2(new_n296), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n247), .B2(new_n296), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n755), .A2(new_n757), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n757), .A2(new_n798), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n752), .B1(new_n756), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n701), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n699), .A2(new_n700), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n809), .B1(new_n812), .B2(new_n752), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT97), .ZN(G396));
  INV_X1    g0614(.A(new_n752), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n446), .A2(new_n694), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n448), .A2(new_n450), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n448), .A2(new_n450), .A3(KEYINPUT99), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n695), .B(new_n821), .C1(new_n681), .C2(new_n685), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n686), .A2(new_n694), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n656), .A2(new_n694), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n819), .A2(new_n824), .A3(new_n820), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n815), .B1(new_n826), .B2(new_n741), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n741), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n757), .A2(new_n753), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT98), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n815), .B1(G77), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n760), .A2(new_n832), .B1(new_n778), .B2(new_n556), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n773), .A2(new_n834), .B1(new_n776), .B2(new_n525), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(new_n770), .C2(G107), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n471), .B1(new_n783), .B2(new_n521), .ZN(new_n837));
  INV_X1    g0637(.A(new_n788), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(G294), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n839), .C1(new_n539), .C2(new_n787), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G150), .A2(new_n774), .B1(new_n777), .B2(new_n762), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n787), .C1(new_n843), .C2(new_n788), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT34), .Z(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n783), .A2(new_n227), .B1(new_n760), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n263), .B1(new_n778), .B2(new_n228), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n202), .B2(new_n769), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n831), .B1(new_n851), .B2(new_n757), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n825), .B2(new_n754), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n828), .A2(new_n853), .ZN(G384));
  NOR2_X1   g0654(.A1(new_n746), .A2(new_n307), .ZN(new_n855));
  INV_X1    g0655(.A(new_n692), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n655), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n448), .A2(new_n694), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n822), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n344), .A2(new_n695), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n384), .A2(new_n387), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(G169), .B1(new_n363), .B2(new_n376), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT14), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n387), .A2(new_n866), .A3(new_n380), .A4(new_n377), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT102), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n862), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n868), .B1(new_n867), .B2(new_n862), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n453), .B(new_n465), .C1(new_n510), .C2(new_n496), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n488), .A2(new_n489), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n513), .B1(new_n454), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT103), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n454), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n505), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n498), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n856), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n498), .B1(new_n511), .B2(new_n692), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n511), .A2(new_n886), .A3(new_n513), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n501), .A2(new_n505), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT37), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n884), .A2(KEYINPUT37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n651), .A2(new_n652), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n498), .A2(new_n499), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT17), .B1(new_n511), .B2(new_n466), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n874), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n883), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n500), .B2(new_n515), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n888), .A2(new_n890), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n498), .A2(new_n881), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n898), .B1(new_n902), .B2(KEYINPUT103), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n903), .B2(new_n882), .ZN(new_n904));
  OAI211_X1 g0704(.A(KEYINPUT38), .B(new_n899), .C1(new_n900), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n857), .B1(new_n873), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n653), .A2(new_n895), .A3(new_n654), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n501), .A2(new_n856), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n888), .A2(new_n890), .ZN(new_n913));
  INV_X1    g0713(.A(new_n889), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n914), .B2(new_n885), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n891), .A2(new_n874), .A3(new_n896), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n908), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n384), .A2(new_n694), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n897), .A2(new_n905), .A3(KEYINPUT39), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n907), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n517), .B1(new_n717), .B2(new_n723), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n664), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n736), .A2(new_n737), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n725), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n825), .C1(new_n870), .C2(new_n871), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT40), .B1(new_n906), .B2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n909), .A2(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n905), .B1(new_n933), .B2(KEYINPUT38), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n932), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n517), .A2(new_n929), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n700), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n855), .B1(new_n927), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n927), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n943));
  OAI211_X1 g0743(.A(G116), .B(new_n226), .C1(new_n625), .C2(KEYINPUT35), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT100), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  XNOR2_X1  g0747(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n475), .A2(G77), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n243), .B1(new_n230), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(G1), .A3(new_n219), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n942), .A2(new_n949), .A3(new_n952), .ZN(G367));
  NOR2_X1   g0753(.A1(new_n803), .A2(new_n241), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n807), .B1(new_n221), .B2(new_n440), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n815), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n778), .A2(new_n521), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n773), .A2(new_n292), .B1(new_n776), .B2(new_n834), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(G107), .C2(new_n784), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n471), .B1(new_n760), .B2(new_n960), .C1(new_n787), .C2(new_n832), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G303), .B2(new_n838), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n769), .B2(new_n525), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n959), .A2(new_n962), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n471), .B1(new_n784), .B2(G68), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n787), .B2(new_n843), .C1(new_n393), .C2(new_n788), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n774), .A2(new_n762), .B1(new_n761), .B2(G137), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n778), .A2(new_n335), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G50), .B2(new_n777), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(new_n227), .C2(new_n769), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n966), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT108), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT47), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n956), .B1(new_n975), .B2(new_n757), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n562), .A2(new_n582), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n694), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n673), .A2(new_n676), .A3(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(new_n676), .C2(new_n978), .ZN(new_n982));
  INV_X1    g0782(.A(new_n755), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n634), .B(new_n646), .C1(new_n640), .C2(new_n695), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n634), .B2(new_n695), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n710), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n710), .A2(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n707), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n709), .A2(new_n329), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n705), .B2(new_n709), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n701), .B(new_n994), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n742), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n743), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n712), .B(KEYINPUT41), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n750), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n986), .B(KEYINPUT107), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n328), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n694), .B1(new_n1003), .B2(new_n634), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n986), .A2(new_n329), .A3(new_n709), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT42), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1001), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT106), .Z(new_n1009));
  XNOR2_X1  g0809(.A(new_n1007), .B(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1002), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n707), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1010), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n984), .B1(new_n1000), .B2(new_n1013), .ZN(G387));
  NOR2_X1   g0814(.A1(new_n996), .A2(new_n745), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n995), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n743), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n783), .A2(new_n440), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n773), .A2(new_n392), .B1(new_n776), .B2(new_n228), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G150), .C2(new_n761), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n787), .A2(new_n477), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT109), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n770), .A2(G77), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n471), .B(new_n957), .C1(new_n838), .C2(G50), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n263), .B1(new_n779), .B2(G116), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n769), .A2(new_n292), .B1(new_n834), .B2(new_n783), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n774), .B1(new_n777), .B2(G303), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n960), .B2(new_n788), .C1(new_n792), .C2(new_n787), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1026), .B1(new_n791), .B2(new_n760), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n757), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n238), .A2(new_n296), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(new_n802), .B1(new_n713), .B2(new_n799), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT50), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n438), .B2(new_n202), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n392), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n296), .B1(new_n228), .B2(new_n335), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n713), .A4(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1039), .A2(new_n1044), .B1(G107), .B2(new_n221), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n752), .B1(new_n1045), .B2(new_n807), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1037), .B(new_n1046), .C1(new_n705), .C2(new_n983), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1017), .B(new_n1047), .C1(new_n747), .C2(new_n995), .ZN(G393));
  AOI21_X1  g0848(.A(new_n745), .B1(new_n992), .B2(new_n996), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n996), .B2(new_n992), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT111), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n1011), .A2(new_n755), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n807), .B1(new_n221), .B2(new_n521), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n802), .B2(new_n250), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n774), .A2(G303), .B1(new_n761), .B2(G322), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n525), .B2(new_n783), .C1(new_n292), .C2(new_n776), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n263), .B(new_n1056), .C1(G107), .C2(new_n779), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n834), .B2(new_n769), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n832), .A2(new_n788), .B1(new_n787), .B2(new_n960), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  OAI22_X1  g0860(.A1(new_n393), .A2(new_n787), .B1(new_n788), .B2(new_n477), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  AOI22_X1  g0862(.A1(new_n774), .A2(G50), .B1(new_n761), .B2(G143), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n784), .A2(G77), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n392), .C2(new_n776), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n471), .B(new_n1065), .C1(G87), .C2(new_n779), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n228), .B2(new_n769), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1058), .A2(new_n1060), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n752), .B(new_n1054), .C1(new_n1068), .C2(new_n757), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT110), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n992), .A2(new_n750), .B1(new_n1052), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1051), .A2(new_n1071), .ZN(G390));
  NAND2_X1  g0872(.A1(new_n919), .A2(new_n922), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n871), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n864), .A3(new_n869), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n921), .B1(new_n860), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n821), .B(new_n695), .C1(new_n685), .C2(new_n720), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1075), .B1(new_n1080), .B2(new_n858), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n920), .B(KEYINPUT112), .Z(new_n1082));
  NAND3_X1  g0882(.A1(new_n934), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1075), .A2(G330), .A3(new_n740), .A4(new_n825), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1078), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n700), .B1(new_n725), .B2(new_n928), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1075), .A2(new_n825), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1076), .B1(new_n919), .B2(new_n922), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1083), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n747), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n769), .A2(new_n393), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  INV_X1    g0895(.A(G128), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n263), .B1(new_n773), .B2(new_n842), .C1(new_n1096), .C2(new_n787), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G132), .B2(new_n838), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n778), .A2(new_n202), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n776), .A2(new_n1100), .B1(new_n783), .B2(new_n477), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G125), .C2(new_n761), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n771), .A2(new_n471), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT114), .Z(new_n1105));
  OAI221_X1 g0905(.A(new_n1064), .B1(new_n228), .B2(new_n778), .C1(new_n788), .C2(new_n525), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n787), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(G283), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G107), .A2(new_n774), .B1(new_n777), .B2(G97), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n292), .C2(new_n760), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1103), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n757), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n815), .B1(new_n438), .B2(new_n830), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(new_n1073), .C2(new_n753), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1093), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n517), .A2(new_n1086), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n925), .A2(new_n1116), .A3(new_n664), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n740), .A2(G330), .A3(new_n825), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n872), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT113), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT113), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1118), .A2(new_n1121), .A3(new_n872), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1087), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n860), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1079), .A2(new_n859), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1086), .A2(new_n825), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n872), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1084), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1117), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1092), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1085), .A2(new_n1129), .A3(new_n1091), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n712), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1115), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT115), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT115), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1115), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G378));
  OAI21_X1  g0939(.A(new_n936), .B1(new_n917), .B2(new_n918), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(G330), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n932), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n906), .A2(new_n931), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n935), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT117), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n700), .B1(new_n934), .B2(new_n936), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n660), .A2(new_n427), .A3(new_n662), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n424), .A2(new_n692), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1152), .B(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1142), .A2(new_n1147), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1153), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1159), .A2(new_n1145), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n924), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n924), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n750), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n263), .A2(G41), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(G33), .A2(G41), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT116), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1166), .A2(new_n1168), .A3(G50), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n778), .A2(new_n227), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n773), .A2(new_n521), .B1(new_n776), .B2(new_n440), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G283), .C2(new_n761), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1166), .B1(new_n783), .B2(new_n228), .C1(new_n788), .C2(new_n254), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G116), .B2(new_n1107), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1023), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1169), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n773), .A2(new_n846), .B1(new_n776), .B2(new_n842), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G150), .B2(new_n784), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G125), .A2(new_n1107), .B1(new_n838), .B2(G128), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n769), .C2(new_n1100), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n779), .A2(new_n762), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n761), .A2(G124), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1168), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n757), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n830), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n752), .B1(new_n202), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(new_n1155), .C2(new_n754), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1156), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1163), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1117), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1132), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1162), .A2(new_n1197), .A3(KEYINPUT57), .A4(new_n1164), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n712), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1192), .B1(new_n1198), .B2(new_n1200), .ZN(G375));
  NAND3_X1  g1001(.A1(new_n1124), .A2(new_n1117), .A3(new_n1128), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT118), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1128), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1123), .B2(new_n860), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT118), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1117), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1130), .A3(new_n999), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n872), .A2(new_n753), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n815), .B1(G68), .B2(new_n830), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1107), .A2(G132), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT121), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n770), .A2(G159), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n776), .A2(new_n393), .B1(new_n783), .B2(new_n202), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n773), .A2(new_n1100), .B1(new_n760), .B2(new_n1096), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n471), .B(new_n1170), .C1(new_n838), .C2(G137), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1213), .A2(new_n1214), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n773), .A2(new_n525), .B1(new_n776), .B2(new_n254), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT119), .Z(new_n1221));
  NOR2_X1   g1021(.A1(new_n760), .A2(new_n539), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1222), .B(new_n1018), .C1(G294), .C2(new_n1107), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(new_n834), .C2(new_n788), .ZN(new_n1224));
  OR3_X1    g1024(.A1(new_n970), .A2(KEYINPUT120), .A3(new_n263), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT120), .B1(new_n970), .B2(new_n263), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n521), .C2(new_n769), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1219), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1211), .B1(new_n1228), .B2(new_n757), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1209), .A2(new_n750), .B1(new_n1210), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1208), .A2(new_n1230), .ZN(G381));
  OR2_X1    g1031(.A1(G393), .A2(G396), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(G390), .A2(G384), .A3(G387), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1134), .ZN(new_n1234));
  INV_X1    g1034(.A(G375), .ZN(new_n1235));
  INV_X1    g1035(.A(G381), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(G407));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(G343), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1234), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(G213), .A3(new_n1240), .ZN(G409));
  NAND2_X1  g1041(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1242));
  XOR2_X1   g1042(.A(G393), .B(G396), .Z(new_n1243));
  MUX2_X1   g1043(.A(new_n1242), .B(G387), .S(new_n1243), .Z(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(G390), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1205), .B2(new_n1117), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1203), .A2(new_n1247), .A3(new_n1207), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1202), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n745), .B1(new_n1249), .B2(KEYINPUT60), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1250), .A3(KEYINPUT123), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G384), .B1(new_n1255), .B2(new_n1230), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1248), .A2(new_n1250), .A3(KEYINPUT123), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT123), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G384), .B(new_n1230), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1239), .A2(G2897), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1162), .A2(new_n1197), .A3(new_n999), .A4(new_n1164), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1165), .A3(new_n1191), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1234), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(G375), .B2(new_n1138), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1239), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1263), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1245), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1267), .A2(new_n1268), .A3(new_n1261), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1267), .A2(KEYINPUT124), .A3(new_n1268), .A4(new_n1261), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1272), .B(new_n1278), .C1(new_n1276), .C2(new_n1273), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1275), .A2(KEYINPUT126), .A3(new_n1280), .A4(new_n1277), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1269), .A2(KEYINPUT62), .A3(new_n1261), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1275), .A2(new_n1280), .A3(new_n1277), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1271), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1244), .B(G390), .Z(new_n1288));
  OAI21_X1  g1088(.A(new_n1279), .B1(new_n1287), .B2(new_n1288), .ZN(G405));
  NOR2_X1   g1089(.A1(new_n1261), .A2(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1245), .B1(KEYINPUT127), .B2(new_n1261), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1261), .A2(KEYINPUT127), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1235), .A2(G378), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1234), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1297), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1291), .A2(new_n1292), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(G402));
endmodule


