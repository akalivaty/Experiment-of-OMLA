//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n441, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1260, new_n1261, new_n1262;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT70), .B1(new_n462), .B2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT69), .B1(new_n462), .B2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n460), .A3(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n470), .A2(G137), .A3(new_n471), .A4(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n460), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n467), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  INV_X1    g055(.A(KEYINPUT73), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n463), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n475), .A2(new_n471), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n484), .B1(new_n489), .B2(G136), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n470), .A2(G2105), .A3(new_n475), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n481), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n490), .A2(new_n493), .A3(new_n481), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  NOR4_X1   g075(.A1(new_n464), .A2(KEYINPUT4), .A3(new_n499), .A4(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n470), .A2(G126), .A3(G2105), .A4(new_n475), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT74), .B(G114), .Z(new_n507));
  OAI211_X1 g082(.A(G2104), .B(new_n506), .C1(new_n507), .C2(new_n471), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n470), .A2(G138), .A3(new_n471), .A4(new_n475), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n501), .B1(new_n512), .B2(KEYINPUT4), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT75), .B1(new_n513), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT76), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G62), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n516), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(G88), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(G50), .A3(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n527), .A2(new_n532), .A3(KEYINPUT77), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n534), .B1(new_n526), .B2(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(G166));
  NAND2_X1  g111(.A1(new_n522), .A2(new_n523), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n538));
  INV_X1    g113(.A(G63), .ZN(new_n539));
  NOR4_X1   g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n516), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n522), .A2(new_n523), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n516), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT78), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(G89), .A3(new_n528), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n528), .A2(G543), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT79), .B(G51), .Z(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT80), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n541), .A2(new_n542), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(new_n538), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n541), .A2(KEYINPUT78), .A3(new_n542), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n552), .A2(new_n559), .ZN(G168));
  NAND2_X1  g135(.A1(G77), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G64), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n537), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n541), .A2(G90), .A3(new_n528), .ZN(new_n565));
  XOR2_X1   g140(.A(KEYINPUT81), .B(G52), .Z(new_n566));
  NAND2_X1  g141(.A1(new_n548), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n565), .A2(KEYINPUT82), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT82), .B1(new_n565), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(G301));
  INV_X1    g145(.A(G301), .ZN(G171));
  AOI22_X1  g146(.A1(new_n541), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n516), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n541), .A2(new_n528), .ZN(new_n574));
  INV_X1    g149(.A(G81), .ZN(new_n575));
  INV_X1    g150(.A(new_n548), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT83), .B(G43), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  AND3_X1   g155(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G36), .ZN(G176));
  NAND2_X1  g157(.A1(G1), .A2(G3), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT8), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G188));
  NAND2_X1  g160(.A1(new_n548), .A2(G53), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n541), .A2(new_n528), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n587), .A2(new_n588), .B1(G91), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT84), .B(G65), .Z(new_n591));
  AOI22_X1  g166(.A1(new_n541), .A2(new_n591), .B1(G78), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n516), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G299));
  AND2_X1   g169(.A1(new_n552), .A2(new_n559), .ZN(G286));
  INV_X1    g170(.A(G166), .ZN(G303));
  NAND2_X1  g171(.A1(new_n589), .A2(G87), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n541), .B2(G74), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n548), .A2(G49), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  AOI22_X1  g175(.A1(new_n541), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n516), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n548), .A2(G48), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n574), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G305));
  AOI22_X1  g183(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n516), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n589), .A2(G85), .B1(G47), .B2(new_n548), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n541), .A2(G92), .A3(new_n528), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n576), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n548), .A2(KEYINPUT85), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n537), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n618), .A2(new_n619), .B1(G651), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n613), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n613), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(G868), .B2(new_n628), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(G868), .B2(new_n628), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n489), .B2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n492), .A2(G123), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2446), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G2443), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(G2443), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n652), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n658), .A2(G2443), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n659), .A3(new_n651), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1341), .B(G1348), .Z(new_n666));
  AOI21_X1  g241(.A(KEYINPUT86), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n662), .A2(new_n664), .ZN(new_n670));
  INV_X1    g245(.A(new_n666), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(KEYINPUT86), .A3(new_n666), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(KEYINPUT17), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n677), .A3(new_n678), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n678), .A2(new_n679), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT18), .Z(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2096), .B(G2100), .Z(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n695), .B(new_n704), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n705), .A2(KEYINPUT20), .A3(new_n697), .A4(new_n698), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n700), .A2(new_n703), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G1991), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(G1991), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(G1996), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(G1996), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n694), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(new_n694), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n716), .A3(new_n711), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n714), .A2(new_n717), .A3(new_n719), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(G229));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G24), .ZN(new_n725));
  INV_X1    g300(.A(G290), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  INV_X1    g303(.A(G25), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G29), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(G107), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n489), .B2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n492), .A2(G119), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT91), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n729), .B2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n731), .B1(new_n743), .B2(KEYINPUT90), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT35), .B(G1991), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n728), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(G16), .A2(G23), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G288), .B2(new_n724), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT33), .B(G1976), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G305), .A2(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n724), .A2(G6), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT32), .B(G1981), .Z(new_n754));
  AND3_X1   g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n751), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G22), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G166), .B2(G16), .ZN(new_n759));
  INV_X1    g334(.A(G1971), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n757), .B(KEYINPUT34), .C1(new_n761), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n746), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n744), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n747), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT36), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n747), .A2(new_n767), .A3(new_n772), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n497), .A2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G29), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G35), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT29), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n775), .A2(new_n780), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G2090), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n784));
  INV_X1    g359(.A(G26), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G29), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(G29), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G116), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n489), .B2(G140), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n492), .A2(G128), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n791), .A2(new_n792), .A3(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n787), .B1(new_n797), .B2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n786), .B1(new_n798), .B2(new_n784), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(G2067), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n783), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G2090), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n779), .A2(new_n802), .A3(new_n781), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(G2067), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT96), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT26), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n477), .A2(G105), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n489), .B2(G141), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n492), .A2(G129), .ZN(new_n814));
  AOI21_X1  g389(.A(KEYINPUT97), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n809), .A2(new_n811), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n489), .A2(G141), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  OR2_X1    g397(.A1(G29), .A2(G32), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT27), .B(G1996), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n477), .A2(G103), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT93), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n827), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT25), .ZN(new_n833));
  NAND2_X1  g408(.A1(G115), .A2(G2104), .ZN(new_n834));
  INV_X1    g409(.A(G127), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n464), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G2105), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n830), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G139), .B2(new_n489), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n776), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n776), .A2(G33), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT94), .B(G2072), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n724), .A2(G4), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n615), .A2(new_n623), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(G16), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(G1348), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(G1348), .ZN(new_n851));
  OAI22_X1  g426(.A1(new_n844), .A2(new_n845), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(G5), .A2(G16), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G171), .B2(G16), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(G1961), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(G1961), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n642), .A2(new_n776), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT99), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT99), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n855), .B(new_n856), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n724), .B1(new_n590), .B2(new_n593), .ZN(new_n861));
  INV_X1    g436(.A(G1956), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n724), .A2(G20), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OR3_X1    g440(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n861), .B2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n724), .A2(G19), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n573), .A2(new_n578), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(G16), .ZN(new_n871));
  INV_X1    g446(.A(G1341), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G2084), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT24), .ZN(new_n875));
  INV_X1    g450(.A(G34), .ZN(new_n876));
  AOI21_X1  g451(.A(G29), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n479), .B2(G29), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT30), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(G28), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n776), .B1(new_n882), .B2(G28), .ZN(new_n884));
  AND2_X1   g459(.A1(KEYINPUT31), .A2(G11), .ZN(new_n885));
  NOR2_X1   g460(.A1(KEYINPUT31), .A2(G11), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n880), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(G2084), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n868), .A2(new_n873), .A3(new_n881), .A4(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n852), .A2(new_n860), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n511), .A2(G29), .A3(new_n514), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n776), .A2(G27), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G2078), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(G2078), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n724), .A2(G21), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G286), .B2(G16), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT98), .B(G1966), .Z(new_n900));
  OR2_X1    g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  AOI211_X1 g477(.A(new_n896), .B(new_n897), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n826), .A2(new_n891), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT101), .B1(new_n806), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n826), .A2(new_n891), .A3(new_n903), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  NOR4_X1   g482(.A1(new_n906), .A2(new_n801), .A3(new_n907), .A4(new_n805), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n774), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(G311));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n774), .B(KEYINPUT102), .C1(new_n905), .C2(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G150));
  NOR2_X1   g489(.A1(new_n848), .A2(new_n631), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n548), .A2(G55), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT103), .B(G93), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n574), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n541), .A2(G67), .ZN(new_n921));
  NAND2_X1  g496(.A1(G80), .A2(G543), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n516), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n579), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G860), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n925), .B2(new_n917), .ZN(new_n927));
  OAI21_X1  g502(.A(G860), .B1(new_n920), .B2(new_n923), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT37), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(G145));
  NAND3_X1  g505(.A1(new_n797), .A2(new_n739), .A3(new_n740), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n741), .A2(new_n795), .A3(new_n796), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n492), .A2(G130), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n489), .A2(G142), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n471), .A2(G118), .ZN(new_n936));
  OAI21_X1  g511(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n513), .A2(new_n509), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n931), .A2(new_n932), .A3(new_n940), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n495), .B(new_n496), .C1(new_n815), .C2(new_n820), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n642), .B(new_n479), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n813), .A2(KEYINPUT97), .A3(new_n814), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n818), .A2(new_n819), .ZN(new_n947));
  INV_X1    g522(.A(new_n496), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n946), .B(new_n947), .C1(new_n494), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n945), .B1(new_n944), .B2(new_n949), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n942), .B(new_n943), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n949), .ZN(new_n954));
  INV_X1    g529(.A(new_n945), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n931), .A2(new_n932), .A3(new_n940), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n940), .B1(new_n931), .B2(new_n932), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n956), .B(new_n950), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n645), .B(KEYINPUT104), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n839), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n953), .A2(new_n959), .ZN(new_n965));
  INV_X1    g540(.A(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n924), .B2(G868), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n870), .B(new_n924), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n633), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n925), .A2(new_n631), .A3(new_n624), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n624), .A2(G299), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n628), .A2(new_n848), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT105), .Z(new_n979));
  INV_X1    g554(.A(KEYINPUT41), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n975), .A2(KEYINPUT41), .A3(new_n976), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n973), .A2(new_n974), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n983), .B2(new_n985), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n979), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n602), .A2(new_n606), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(G290), .ZN(new_n992));
  XNOR2_X1  g567(.A(G166), .B(G288), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n991), .B(new_n726), .ZN(new_n995));
  INV_X1    g570(.A(new_n993), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n979), .B(new_n1000), .C1(new_n986), .C2(new_n987), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n989), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G868), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n999), .B1(new_n989), .B2(new_n1001), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n971), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n989), .A2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n998), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(new_n970), .A3(G868), .A4(new_n1002), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(G295));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1008), .ZN(G331));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n1011));
  INV_X1    g586(.A(new_n569), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n565), .A2(KEYINPUT82), .A3(new_n567), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n1014), .B2(new_n564), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1011), .B(new_n564), .C1(new_n568), .C2(new_n569), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G168), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G301), .A2(KEYINPUT109), .ZN(new_n1019));
  NAND3_X1  g594(.A1(G286), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1020), .A3(new_n925), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1018), .A2(new_n1020), .A3(KEYINPUT110), .A4(new_n925), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1026), .A2(new_n972), .B1(new_n976), .B2(new_n975), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n972), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1021), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1025), .A2(new_n1027), .B1(new_n1029), .B2(new_n983), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n998), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G37), .B1(new_n1030), .B2(new_n998), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT43), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1025), .A2(new_n1028), .B1(new_n981), .B2(new_n982), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1027), .A2(new_n1021), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n999), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1033), .A2(new_n1037), .A3(KEYINPUT43), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT44), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1029), .A2(new_n983), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n998), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n963), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT43), .B1(new_n1043), .B2(new_n1031), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1033), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1039), .B1(new_n1048), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g624(.A(G1384), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n513), .B2(new_n509), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n467), .A2(new_n476), .A3(G40), .A4(new_n478), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n797), .A2(G2067), .ZN(new_n1057));
  INV_X1    g632(.A(G2067), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n795), .A2(new_n1058), .A3(new_n796), .ZN(new_n1059));
  INV_X1    g634(.A(G1996), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1057), .B(new_n1059), .C1(new_n821), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT111), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1061), .A2(new_n1055), .B1(new_n1063), .B2(new_n821), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(new_n768), .A3(new_n739), .A4(new_n740), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1056), .B1(new_n1065), .B2(new_n1059), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n741), .B(new_n746), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1056), .B1(new_n1067), .B2(KEYINPUT112), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(KEYINPUT112), .B2(new_n1067), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1056), .A2(G1986), .A3(G290), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1070), .B(KEYINPUT48), .Z(new_n1071));
  AND3_X1   g646(.A1(new_n1069), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1063), .B(KEYINPUT46), .Z(new_n1073));
  AND3_X1   g648(.A1(new_n1057), .A2(new_n821), .A3(new_n1059), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1056), .B2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1075), .A2(KEYINPUT47), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(KEYINPUT47), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1066), .B(new_n1072), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G288), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G1976), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT52), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT49), .ZN(new_n1086));
  INV_X1    g661(.A(G1981), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n603), .B2(new_n607), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n602), .A2(new_n606), .A3(G1981), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n990), .A2(new_n1087), .ZN(new_n1091));
  OAI21_X1  g666(.A(G1981), .B1(new_n602), .B2(new_n606), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT49), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1081), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1976), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(G288), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1081), .A2(new_n1083), .A3(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1085), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n511), .A2(new_n1050), .A3(new_n514), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT50), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n1050), .C1(new_n513), .C2(new_n509), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1054), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1103), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1052), .B2(new_n1099), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1106), .A2(G2090), .B1(new_n1108), .B2(G1971), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n533), .A2(G8), .A3(new_n535), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1111), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n533), .A2(new_n535), .A3(G8), .A4(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1109), .A2(new_n1118), .A3(G8), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n511), .A2(new_n514), .A3(new_n1101), .A4(new_n1050), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1054), .B1(new_n1051), .B2(KEYINPUT50), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT116), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1124), .A3(new_n1121), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n802), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1099), .A2(new_n1052), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1107), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n760), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1080), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1098), .B(new_n1119), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1104), .B1(new_n1099), .B2(KEYINPUT50), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT45), .A4(new_n1050), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(new_n1103), .A3(new_n1053), .ZN(new_n1136));
  INV_X1    g711(.A(new_n900), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n874), .A2(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1138), .A2(new_n1080), .A3(G286), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT117), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1119), .A2(new_n1098), .ZN(new_n1143));
  AOI21_X1  g718(.A(G2090), .B1(new_n1122), .B2(KEYINPUT116), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1144), .A2(new_n1125), .B1(new_n760), .B2(new_n1129), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1115), .B(new_n1112), .C1(new_n1145), .C2(new_n1080), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .A4(new_n1139), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1141), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1109), .A2(G8), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1132), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(KEYINPUT63), .A3(new_n1143), .A4(new_n1139), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1098), .A2(G8), .A3(new_n1109), .A4(new_n1118), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1094), .A2(new_n1095), .A3(new_n1082), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1081), .B1(new_n1157), .B2(new_n1089), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G286), .A2(G8), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1134), .A2(new_n874), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1080), .B1(new_n1138), .B2(G168), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(KEYINPUT51), .B(new_n1161), .C1(new_n1138), .C2(new_n1080), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT123), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1166), .B(G8), .C1(new_n1170), .C2(G286), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1164), .ZN(new_n1172));
  AND4_X1   g747(.A1(KEYINPUT123), .A2(new_n1171), .A3(new_n1168), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT62), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT53), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1129), .B2(G2078), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1134), .A2(G1961), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1175), .B(G2078), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(new_n1103), .A3(new_n1135), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(G301), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1167), .A2(KEYINPUT123), .A3(new_n1168), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1171), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1174), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT56), .B(G2072), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1108), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1122), .A2(new_n862), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G299), .B(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1079), .A2(new_n1058), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT120), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1134), .A2(G1348), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n848), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1195), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1190), .A2(new_n1194), .A3(new_n1204), .A4(new_n1191), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(KEYINPUT61), .ZN(new_n1206));
  AOI21_X1  g781(.A(KEYINPUT122), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1207));
  OR2_X1    g782(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1129), .A2(G1996), .ZN(new_n1210));
  XNOR2_X1  g785(.A(KEYINPUT58), .B(G1341), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1079), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n579), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1199), .A2(new_n1216), .A3(new_n1201), .A4(new_n1217), .ZN(new_n1218));
  OAI211_X1 g793(.A(KEYINPUT60), .B(new_n624), .C1(new_n1198), .C2(new_n1200), .ZN(new_n1219));
  OAI211_X1 g794(.A(KEYINPUT59), .B(new_n579), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1215), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1203), .B1(new_n1209), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n476), .A2(new_n478), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n1224));
  OAI211_X1 g799(.A(G40), .B(new_n467), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1225), .B1(new_n1224), .B2(new_n1223), .ZN(new_n1226));
  OAI211_X1 g801(.A(new_n1178), .B(new_n1226), .C1(new_n1052), .C2(new_n1051), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1176), .A2(new_n1177), .A3(G301), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1228), .B1(new_n1180), .B2(G301), .ZN(new_n1229));
  XNOR2_X1  g804(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1180), .A2(G301), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT54), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1176), .A2(new_n1177), .A3(new_n1227), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1232), .B1(new_n1233), .B2(G171), .ZN(new_n1234));
  AOI22_X1  g809(.A1(new_n1229), .A2(new_n1230), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g810(.A(new_n1222), .B(new_n1235), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1188), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(new_n1133), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1160), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g814(.A(G290), .B(G1986), .Z(new_n1240));
  OAI211_X1 g815(.A(new_n1069), .B(new_n1064), .C1(new_n1056), .C2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g816(.A(new_n1241), .B(KEYINPUT113), .Z(new_n1242));
  OAI21_X1  g817(.A(new_n1078), .B1(new_n1239), .B2(new_n1242), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g818(.A1(new_n691), .A2(G319), .A3(new_n692), .ZN(new_n1245));
  NAND4_X1  g819(.A1(new_n674), .A2(new_n721), .A3(new_n1245), .A4(new_n722), .ZN(new_n1246));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g822(.A1(new_n691), .A2(G319), .A3(new_n692), .ZN(new_n1249));
  OAI21_X1  g823(.A(G14), .B1(new_n665), .B2(new_n666), .ZN(new_n1250));
  NOR2_X1   g824(.A1(new_n1250), .A2(new_n667), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n1249), .B1(new_n1251), .B2(new_n673), .ZN(new_n1252));
  NAND4_X1  g826(.A1(new_n1252), .A2(KEYINPUT126), .A3(new_n722), .A4(new_n721), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g828(.A(new_n1254), .B1(new_n964), .B2(new_n967), .ZN(new_n1255));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1256));
  AND3_X1   g830(.A1(new_n1255), .A2(new_n1047), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g831(.A(new_n1256), .B1(new_n1255), .B2(new_n1047), .ZN(new_n1258));
  NOR2_X1   g832(.A1(new_n1257), .A2(new_n1258), .ZN(G308));
  NAND2_X1  g833(.A1(new_n1255), .A2(new_n1047), .ZN(new_n1260));
  NAND2_X1  g834(.A1(new_n1260), .A2(KEYINPUT127), .ZN(new_n1261));
  NAND3_X1  g835(.A1(new_n1255), .A2(new_n1047), .A3(new_n1256), .ZN(new_n1262));
  NAND2_X1  g836(.A1(new_n1261), .A2(new_n1262), .ZN(G225));
endmodule


