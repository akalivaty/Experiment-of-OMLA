//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G101), .ZN(new_n197));
  AOI21_X1  g011(.A(G101), .B1(new_n189), .B2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n190), .A2(new_n198), .A3(new_n193), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n195), .B2(G101), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n188), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n201), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n190), .A2(new_n198), .A3(new_n193), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT4), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT77), .A4(new_n197), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G116), .B(G119), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n195), .A2(new_n205), .A3(G101), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G119), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n209), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(new_n218), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n210), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n189), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n192), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n229), .A2(new_n199), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n229), .B2(new_n199), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n214), .B1(new_n202), .B2(new_n207), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .A3(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n248), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n260), .A3(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n256), .B1(G125), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT85), .B(G224), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n265), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n256), .B(new_n267), .C1(G125), .C2(new_n262), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n216), .A2(new_n235), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n236), .A2(KEYINPUT6), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT84), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT84), .B(new_n271), .C1(new_n239), .C2(new_n234), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n241), .B(new_n269), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G101), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n192), .A2(G104), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n194), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n204), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT79), .B1(new_n204), .B2(new_n278), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n229), .A2(new_n199), .A3(new_n230), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n209), .A2(KEYINPUT5), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n224), .B1(new_n221), .B2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n226), .A2(new_n280), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n236), .B(KEYINPUT8), .Z(new_n287));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n288));
  OAI22_X1  g102(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n268), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n267), .A2(KEYINPUT7), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n263), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT86), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n262), .A2(G125), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n248), .A2(new_n251), .B1(new_n249), .B2(new_n253), .ZN(new_n295));
  INV_X1    g109(.A(G125), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n293), .B(new_n290), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n289), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n299), .B2(new_n237), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n275), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n275), .B2(new_n300), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n187), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n275), .A2(new_n300), .ZN(new_n307));
  INV_X1    g121(.A(new_n301), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n275), .A2(new_n300), .A3(new_n301), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT87), .A3(new_n187), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G221), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G113), .B(G122), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(new_n189), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(new_n246), .ZN(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n324), .A2(G143), .A3(G214), .ZN(new_n325));
  AOI21_X1  g139(.A(G143), .B1(new_n324), .B2(G214), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT18), .B(G131), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(G214), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n243), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(G143), .A3(G214), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n296), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT16), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n296), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G146), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(G146), .B1(new_n338), .B2(new_n339), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT17), .B(G131), .C1(new_n325), .C2(new_n326), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n334), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n339), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n246), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(new_n344), .A3(new_n334), .A4(new_n340), .ZN(new_n348));
  OAI21_X1  g162(.A(G131), .B1(new_n325), .B2(new_n326), .ZN(new_n349));
  INV_X1    g163(.A(G131), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n329), .A2(new_n350), .A3(new_n330), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT17), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n321), .B(new_n333), .C1(new_n345), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n351), .ZN(new_n356));
  AND2_X1   g170(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n322), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n322), .B2(new_n358), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n356), .B(new_n340), .C1(new_n360), .C2(G146), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n333), .ZN(new_n362));
  INV_X1    g176(.A(new_n321), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT90), .B1(new_n355), .B2(new_n364), .ZN(new_n369));
  OAI22_X1  g183(.A1(new_n366), .A2(new_n368), .B1(new_n369), .B2(KEYINPUT20), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n368), .B1(new_n355), .B2(new_n364), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n355), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n347), .A2(new_n344), .A3(new_n340), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT89), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n353), .A3(new_n348), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n321), .B1(new_n379), .B2(new_n333), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n317), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n370), .A2(new_n375), .B1(G475), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G953), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n383), .A2(G952), .ZN(new_n384));
  NAND2_X1  g198(.A1(G234), .A2(G237), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(G902), .A3(G953), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT21), .B(G898), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G217), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n315), .A2(new_n393), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n243), .A2(G128), .ZN(new_n396));
  INV_X1    g210(.A(G128), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G134), .ZN(new_n400));
  INV_X1    g214(.A(G134), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G116), .B(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n192), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n219), .A2(KEYINPUT14), .A3(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G107), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(new_n404), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT91), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n404), .A2(new_n409), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n408), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n406), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n404), .B(new_n192), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n402), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT13), .B1(new_n243), .B2(G128), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n397), .B2(G143), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n243), .A2(KEYINPUT13), .A3(G128), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n401), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n395), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n419), .A2(new_n420), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n416), .B(new_n402), .C1(new_n424), .C2(new_n401), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n414), .A2(new_n411), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(new_n394), .C1(new_n426), .C2(new_n406), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AOI211_X1 g246(.A(G902), .B(new_n430), .C1(new_n423), .C2(new_n427), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n382), .A2(new_n392), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT78), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n261), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n253), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n258), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n253), .A2(KEYINPUT78), .A3(new_n260), .A4(G128), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT10), .B1(new_n442), .B2(new_n279), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n262), .A2(KEYINPUT10), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT80), .B1(new_n233), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT10), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n259), .B2(new_n261), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n447), .B(new_n448), .C1(new_n232), .C2(new_n231), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n443), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT69), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n295), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n213), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n208), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT11), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n401), .B2(G137), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT11), .A3(G134), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n401), .A2(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n457), .A2(new_n459), .A3(new_n350), .A4(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(KEYINPUT66), .A3(G131), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(KEYINPUT70), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n450), .A2(new_n455), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  INV_X1    g287(.A(G227), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n473), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n465), .A2(KEYINPUT70), .A3(new_n466), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT70), .B1(new_n465), .B2(new_n466), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n442), .A2(new_n279), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n283), .B2(new_n262), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT12), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n465), .A2(KEYINPUT12), .A3(new_n466), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n450), .A2(new_n455), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT82), .B1(new_n488), .B2(new_n481), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n490), .B(new_n471), .C1(new_n450), .C2(new_n455), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n472), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n492), .B2(new_n476), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n493), .A2(G469), .A3(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n472), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n476), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n472), .A2(KEYINPUT81), .A3(new_n477), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n489), .B2(new_n491), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT81), .B1(new_n472), .B2(new_n477), .ZN(new_n499));
  OAI211_X1 g313(.A(G469), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G469), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n317), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n319), .B(new_n436), .C1(new_n494), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n295), .B(KEYINPUT69), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n469), .A2(new_n507), .A3(new_n470), .ZN(new_n508));
  INV_X1    g322(.A(new_n460), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n401), .A2(G137), .ZN(new_n510));
  OAI21_X1  g324(.A(G131), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n464), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n261), .B2(new_n259), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n508), .A2(new_n211), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT72), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n211), .B1(new_n508), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT28), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n211), .A3(new_n514), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n324), .A2(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT27), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(G101), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT29), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n317), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n530));
  NAND3_X1  g344(.A1(new_n465), .A2(new_n295), .A3(new_n466), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n465), .A2(KEYINPUT67), .A3(new_n295), .A4(new_n466), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n512), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n511), .A2(KEYINPUT68), .A3(new_n464), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n262), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n212), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n530), .B1(new_n519), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n513), .B1(new_n481), .B2(new_n507), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT28), .B1(new_n542), .B2(new_n211), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n527), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n508), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n547), .A3(new_n212), .ZN(new_n548));
  INV_X1    g362(.A(new_n527), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n519), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT29), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G472), .B1(new_n529), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n545), .A2(new_n547), .A3(new_n212), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n519), .A2(new_n527), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT31), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n549), .B1(new_n541), .B2(new_n543), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n548), .A2(new_n557), .A3(new_n527), .A4(new_n519), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n552), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n397), .A2(KEYINPUT23), .A3(G119), .ZN(new_n565));
  INV_X1    g379(.A(G119), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n397), .A2(G119), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n565), .B(new_n567), .C1(new_n569), .C2(KEYINPUT23), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n567), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  OAI22_X1  g386(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n322), .A2(new_n246), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n340), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(G110), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT73), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT73), .B1(new_n571), .B2(new_n572), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n575), .B1(new_n579), .B2(new_n343), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT22), .B(G137), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n383), .A2(G221), .A3(G234), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n317), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(KEYINPUT25), .A3(new_n317), .A4(new_n586), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(KEYINPUT74), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n393), .B1(G234), .B2(new_n317), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT74), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(new_n593), .A3(new_n588), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n592), .A2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n586), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n564), .A2(KEYINPUT75), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT75), .B1(new_n564), .B2(new_n599), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n313), .B(new_n506), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  INV_X1    g417(.A(new_n443), .ZN(new_n604));
  INV_X1    g418(.A(new_n449), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n448), .B1(new_n283), .B2(new_n447), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n451), .A2(new_n213), .A3(new_n453), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n202), .B2(new_n207), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n481), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n490), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n488), .A2(KEYINPUT82), .A3(new_n481), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n477), .B1(new_n613), .B2(new_n472), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n501), .B(new_n317), .C1(new_n614), .C2(new_n487), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n503), .A3(new_n500), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n559), .A2(new_n317), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(G472), .B1(new_n561), .B2(new_n559), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n319), .A3(new_n618), .A4(new_n599), .ZN(new_n619));
  INV_X1    g433(.A(new_n187), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n309), .B2(new_n310), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT33), .B1(new_n394), .B2(KEYINPUT92), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n423), .A2(new_n427), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n423), .B2(new_n427), .ZN(new_n625));
  OAI21_X1  g439(.A(G478), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n429), .A2(new_n317), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n428), .B2(new_n429), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n370), .A2(new_n375), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n381), .A2(G475), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n621), .A2(new_n392), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n619), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT93), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  AND2_X1   g451(.A1(new_n374), .A2(new_n373), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n374), .A2(new_n373), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n631), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n434), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n391), .B(KEYINPUT94), .Z(new_n642));
  NAND3_X1  g456(.A1(new_n621), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n619), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NAND2_X1  g460(.A1(new_n306), .A2(new_n312), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n580), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n596), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n595), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n647), .A2(new_n505), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT37), .B(G110), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  AND3_X1   g469(.A1(new_n564), .A2(new_n319), .A3(new_n616), .ZN(new_n656));
  INV_X1    g470(.A(new_n651), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n389), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n386), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n641), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n304), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  AND2_X1   g478(.A1(new_n500), .A2(new_n503), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n318), .B1(new_n665), .B2(new_n615), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n660), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n559), .A2(new_n561), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT32), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n548), .A2(new_n519), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n527), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n515), .A2(new_n517), .ZN(new_n678));
  AOI21_X1  g492(.A(G902), .B1(new_n678), .B2(new_n549), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n311), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n309), .A2(KEYINPUT38), .A3(new_n310), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n374), .B1(new_n372), .B2(new_n373), .ZN(new_n688));
  AND4_X1   g502(.A1(KEYINPUT90), .A2(new_n365), .A3(new_n373), .A4(new_n367), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n631), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n434), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n187), .A3(new_n691), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n683), .A2(new_n651), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n670), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  INV_X1    g509(.A(KEYINPUT96), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n564), .A2(new_n319), .A3(new_n616), .ZN(new_n697));
  INV_X1    g511(.A(new_n629), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n690), .A2(new_n698), .A3(new_n660), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT95), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT95), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n632), .A2(new_n701), .A3(new_n660), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n621), .A2(new_n651), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n696), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n621), .A2(new_n651), .A3(new_n700), .A4(new_n702), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(KEYINPUT96), .A3(new_n666), .A4(new_n564), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  OAI21_X1  g522(.A(G469), .B1(new_n493), .B2(G902), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n615), .ZN(new_n711));
  OAI211_X1 g525(.A(KEYINPUT97), .B(G469), .C1(new_n493), .C2(G902), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n319), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT98), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n318), .B1(new_n711), .B2(new_n712), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT98), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n564), .A2(new_n599), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n633), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  AND2_X1   g537(.A1(new_n715), .A2(new_n718), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n719), .A2(new_n643), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT99), .B(G116), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G18));
  NOR3_X1   g542(.A1(new_n304), .A2(new_n657), .A3(new_n435), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n716), .A2(new_n564), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NAND3_X1  g545(.A1(new_n621), .A2(new_n690), .A3(new_n691), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n617), .A2(G472), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n523), .A2(new_n549), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n555), .A2(new_n558), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n561), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n736), .A3(new_n599), .ZN(new_n737));
  INV_X1    g551(.A(new_n642), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n732), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n724), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT100), .B(G122), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G24));
  AOI211_X1 g556(.A(new_n304), .B(new_n318), .C1(new_n711), .C2(new_n712), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n736), .A3(new_n651), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT101), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n701), .B1(new_n632), .B2(new_n660), .ZN(new_n746));
  INV_X1    g560(.A(new_n660), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n382), .A2(KEYINPUT95), .A3(new_n629), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n700), .A2(new_n702), .A3(KEYINPUT101), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n744), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n302), .A2(new_n303), .A3(new_n620), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n666), .A2(new_n564), .A3(new_n599), .A4(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n700), .A2(new_n702), .A3(KEYINPUT101), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT101), .B1(new_n700), .B2(new_n702), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n754), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n755), .B(new_n319), .C1(new_n494), .C2(new_n504), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n749), .A2(new_n750), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n598), .B1(new_n674), .B2(new_n552), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR2_X1   g581(.A1(new_n756), .A2(new_n661), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n401), .ZN(G36));
  OAI21_X1  g583(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n501), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n502), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n615), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n319), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n667), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n382), .A2(KEYINPUT43), .A3(new_n698), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT102), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n629), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n626), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n382), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT103), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT103), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n782), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n618), .A2(new_n657), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n755), .B1(new_n794), .B2(KEYINPUT44), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT104), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT104), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n798), .A3(KEYINPUT44), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n795), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n780), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n777), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT47), .B(new_n319), .C1(new_n775), .C2(new_n776), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n755), .A2(new_n598), .A3(new_n700), .A4(new_n702), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n564), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n382), .A2(new_n691), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n738), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n306), .A2(new_n312), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n619), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n811), .B1(new_n653), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n619), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n306), .A2(new_n312), .A3(new_n813), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n652), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n313), .A2(new_n506), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n821), .A3(KEYINPUT108), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n719), .A2(new_n761), .ZN(new_n824));
  INV_X1    g638(.A(new_n661), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n824), .A2(new_n825), .B1(new_n751), .B2(new_n762), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n434), .A2(new_n660), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(new_n640), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n432), .A2(new_n433), .A3(new_n747), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n374), .B(new_n373), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT109), .A4(new_n631), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n651), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n309), .A2(new_n187), .A3(new_n310), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n666), .A2(new_n835), .A3(new_n564), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n666), .A2(new_n835), .A3(KEYINPUT110), .A4(new_n564), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n826), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n632), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n738), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n306), .A2(new_n312), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT107), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT107), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n306), .A2(new_n312), .A3(new_n846), .A4(new_n843), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n817), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n602), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n823), .A2(new_n841), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n715), .B(new_n718), .C1(new_n725), .C2(new_n739), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n721), .A2(new_n851), .A3(new_n766), .A4(new_n730), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n743), .A2(new_n751), .B1(new_n656), .B2(new_n662), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n319), .B1(new_n494), .B2(new_n504), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n732), .A2(new_n854), .A3(new_n747), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n657), .A3(new_n682), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n707), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT52), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(new_n707), .A3(new_n859), .A4(new_n856), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n850), .A2(new_n852), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n851), .A2(new_n766), .A3(new_n721), .A4(new_n730), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n816), .A2(new_n822), .A3(new_n602), .A4(new_n848), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n841), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n858), .A2(new_n860), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n737), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n789), .A2(new_n791), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n387), .B(new_n870), .C1(new_n871), .C2(new_n782), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n834), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT106), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n713), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n318), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(KEYINPUT113), .A3(new_n318), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n873), .B1(new_n880), .B2(new_n806), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n714), .A2(new_n834), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n599), .A2(new_n387), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n382), .A2(new_n629), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n882), .A2(new_n683), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n744), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n792), .A2(new_n386), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n892));
  XOR2_X1   g706(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n893));
  AOI21_X1  g707(.A(new_n187), .B1(new_n685), .B2(new_n686), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n716), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(new_n893), .C1(new_n872), .C2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n792), .A2(new_n386), .A3(new_n737), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(KEYINPUT50), .A3(new_n716), .A4(new_n894), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n893), .B1(new_n872), .B2(new_n895), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n891), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT51), .B1(new_n881), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n804), .A2(new_n876), .A3(new_n805), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n873), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n898), .A3(new_n896), .ZN(new_n906));
  INV_X1    g720(.A(new_n891), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT51), .A4(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n882), .A2(new_n632), .A3(new_n683), .A4(new_n884), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n897), .A2(new_n743), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n384), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n882), .A2(new_n889), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n912), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT48), .B1(new_n912), .B2(new_n719), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n903), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n861), .A2(new_n862), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n864), .A2(new_n862), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT111), .B1(new_n865), .B2(new_n841), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n816), .A2(new_n822), .ZN(new_n921));
  INV_X1    g735(.A(new_n841), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT111), .ZN(new_n923));
  INV_X1    g737(.A(new_n849), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n867), .A2(new_n919), .A3(new_n920), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n869), .A2(new_n917), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT116), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n875), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT49), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(KEYINPUT49), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n698), .A2(new_n187), .A3(new_n319), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n598), .A2(new_n936), .A3(new_n690), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT105), .Z(new_n938));
  AND3_X1   g752(.A1(new_n938), .A2(new_n683), .A3(new_n687), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n934), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT117), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT117), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n932), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(G75));
  NOR2_X1   g759(.A1(new_n383), .A2(G952), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n241), .B1(new_n272), .B2(new_n274), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n269), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n918), .A2(new_n926), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(G902), .ZN(new_n951));
  INV_X1    g765(.A(G210), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT119), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(KEYINPUT118), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n949), .A2(KEYINPUT119), .ZN(new_n958));
  OAI221_X1 g772(.A(new_n955), .B1(KEYINPUT118), .B2(new_n958), .C1(new_n951), .C2(new_n952), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n946), .B1(new_n957), .B2(new_n959), .ZN(G51));
  XNOR2_X1  g774(.A(new_n502), .B(KEYINPUT57), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n918), .A2(new_n926), .A3(new_n927), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n927), .B1(new_n918), .B2(new_n926), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT120), .ZN(new_n965));
  INV_X1    g779(.A(new_n493), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n967), .B(new_n961), .C1(new_n962), .C2(new_n963), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n951), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n772), .A3(new_n773), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n946), .B1(new_n969), .B2(new_n971), .ZN(G54));
  NAND2_X1  g786(.A1(KEYINPUT58), .A2(G475), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n366), .B1(new_n951), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n946), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n951), .A2(new_n366), .A3(new_n973), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G60));
  NOR2_X1   g792(.A1(new_n962), .A2(new_n963), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n624), .A2(new_n625), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n627), .B(KEYINPUT59), .Z(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n975), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n869), .A2(new_n928), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n984), .B2(new_n981), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n918), .B2(new_n926), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n585), .A2(new_n586), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n946), .B1(new_n989), .B2(new_n649), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT121), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT61), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  AOI211_X1 g811(.A(KEYINPUT121), .B(new_n997), .C1(new_n992), .C2(new_n993), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(G66));
  OAI21_X1  g813(.A(G953), .B1(new_n264), .B2(new_n390), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n851), .A2(new_n721), .A3(new_n730), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n865), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n947), .B1(G898), .B2(new_n383), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  AOI22_X1  g819(.A1(new_n780), .A2(new_n800), .B1(new_n806), .B2(new_n808), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n842), .A2(new_n812), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(KEYINPUT122), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n755), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n1009), .B(new_n668), .C1(KEYINPUT122), .C2(new_n1007), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n601), .B2(new_n600), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n694), .A2(new_n1012), .A3(new_n707), .A4(new_n853), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n694), .A2(new_n707), .A3(new_n853), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1006), .A2(new_n1011), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n1016), .A2(new_n383), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n545), .A2(new_n547), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(new_n360), .ZN(new_n1019));
  OR3_X1    g833(.A1(new_n1017), .A2(KEYINPUT123), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G900), .A2(G953), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n853), .A2(new_n707), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n719), .A2(new_n732), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n780), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n768), .B1(new_n760), .B2(new_n765), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1006), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1019), .B(new_n1021), .C1(new_n1026), .C2(G953), .ZN(new_n1027));
  OAI21_X1  g841(.A(KEYINPUT123), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1020), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(G953), .B1(new_n474), .B2(new_n658), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT124), .Z(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1020), .A2(new_n1031), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(G72));
  XOR2_X1   g849(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1036));
  NOR2_X1   g850(.A1(new_n675), .A2(new_n317), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1002), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1038), .B1(new_n1016), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1040), .A2(new_n527), .A3(new_n676), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT126), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1040), .A2(KEYINPUT126), .A3(new_n527), .A4(new_n676), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n550), .A2(new_n1038), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n677), .B(new_n1045), .C1(new_n863), .C2(new_n868), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1038), .B1(new_n1026), .B2(new_n1039), .ZN(new_n1047));
  INV_X1    g861(.A(new_n550), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n946), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(KEYINPUT127), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1049), .A2(new_n1046), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT127), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1052), .A2(new_n1053), .A3(new_n1044), .A4(new_n1043), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1051), .A2(new_n1054), .ZN(G57));
endmodule


