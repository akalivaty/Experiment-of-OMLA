//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n474), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n474), .A2(new_n469), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n469), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n491), .A2(new_n492), .A3(new_n490), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n493), .A2(new_n494), .B1(new_n484), .B2(G126), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n469), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT6), .B1(new_n504), .B2(KEYINPUT69), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT70), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT69), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(new_n502), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .B1(KEYINPUT69), .B2(new_n507), .ZN(new_n516));
  INV_X1    g091(.A(new_n510), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NOR3_X1   g093(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n505), .A2(new_n513), .A3(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(new_n512), .A2(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n519), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n502), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n504), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n519), .A2(G52), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(G81), .A2(new_n512), .B1(new_n519), .B2(G43), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n504), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g118(.A1(new_n540), .A2(KEYINPUT72), .A3(new_n504), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n500), .A2(new_n553), .A3(new_n501), .ZN(new_n554));
  AND2_X1   g129(.A1(KEYINPUT5), .A2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(KEYINPUT5), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(G91), .B2(new_n512), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n516), .A2(new_n517), .ZN(new_n563));
  AND2_X1   g138(.A1(KEYINPUT73), .A2(G53), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(KEYINPUT9), .A3(G543), .A4(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n509), .A2(G543), .A3(new_n510), .A4(new_n564), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n566), .B1(new_n565), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n537), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n533), .A2(new_n535), .A3(new_n536), .A4(KEYINPUT76), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G301));
  NAND2_X1  g152(.A1(new_n512), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n519), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n582), .A2(new_n583), .A3(new_n504), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n582), .B2(new_n504), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n584), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(G86), .A2(new_n512), .B1(new_n519), .B2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n555), .A2(new_n556), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n504), .B1(new_n596), .B2(KEYINPUT79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(KEYINPUT79), .B2(new_n596), .ZN(new_n598));
  AOI22_X1  g173(.A1(G85), .A2(new_n512), .B1(new_n519), .B2(G47), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n599), .B2(new_n598), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(new_n519), .A2(G54), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n554), .B2(new_n557), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n509), .A2(G92), .A3(new_n502), .A4(new_n510), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n605), .B(new_n609), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n576), .B2(G868), .ZN(G284));
  AOI21_X1  g191(.A(new_n615), .B1(new_n576), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(G286), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n558), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G91), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n620), .A2(new_n504), .B1(new_n621), .B2(new_n511), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n567), .A2(new_n568), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n567), .A2(new_n568), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT74), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n619), .B1(new_n628), .B2(new_n618), .ZN(G297));
  AOI21_X1  g204(.A(new_n619), .B1(new_n628), .B2(new_n618), .ZN(G280));
  INV_X1    g205(.A(new_n614), .ZN(new_n631));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G860), .ZN(G148));
  NOR2_X1   g208(.A1(new_n614), .A2(G559), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT82), .ZN(new_n635));
  MUX2_X1   g210(.A(new_n545), .B(new_n635), .S(G868), .Z(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n482), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n484), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n469), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n482), .A2(G2104), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT13), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n661), .A2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT86), .Z(new_n668));
  AND2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n682), .A2(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  INV_X1    g264(.A(new_n685), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n682), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n695), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G33), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT25), .Z(new_n705));
  INV_X1    g280(.A(G139), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n470), .B2(new_n706), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(new_n469), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT93), .Z(new_n711));
  AOI21_X1  g286(.A(new_n703), .B1(new_n711), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2072), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NOR2_X1   g289(.A1(G171), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G5), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n714), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n716), .A2(new_n717), .B1(new_n719), .B2(G1966), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n719), .A2(G1966), .ZN(new_n722));
  NOR2_X1   g297(.A1(G27), .A2(G29), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G164), .B2(G29), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2078), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT24), .ZN(new_n726));
  INV_X1    g301(.A(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n726), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G160), .B2(new_n702), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n702), .A2(G35), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n488), .B2(G29), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G2090), .ZN(new_n737));
  NOR4_X1   g312(.A1(new_n721), .A2(new_n722), .A3(new_n725), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n714), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT23), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n627), .B2(new_n714), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n702), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n484), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n463), .A2(G105), .ZN(new_n749));
  INV_X1    g324(.A(G141), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n470), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n744), .B1(new_n752), .B2(new_n702), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n702), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n482), .A2(G140), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n484), .A2(G128), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n469), .A2(G116), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n702), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n643), .B2(new_n702), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n755), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n714), .A2(G19), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT92), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n546), .B2(new_n714), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1341), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n736), .A2(G2090), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n716), .B2(new_n717), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n771), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n730), .A2(G2084), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  NOR2_X1   g355(.A1(G4), .A2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT91), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n614), .B2(new_n714), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n738), .A2(new_n743), .A3(new_n778), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT97), .ZN(new_n788));
  NOR2_X1   g363(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n789));
  MUX2_X1   g364(.A(G6), .B(G305), .S(G16), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT32), .B(G1981), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n714), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n714), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n714), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n714), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT33), .B(G1976), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n792), .A2(KEYINPUT34), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n603), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G16), .B2(G24), .ZN(new_n804));
  INV_X1    g379(.A(G1986), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n702), .A2(G25), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n482), .A2(G131), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT89), .Z(new_n810));
  OR2_X1    g385(.A1(new_n469), .A2(G107), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n484), .A2(G119), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n808), .B1(new_n816), .B2(new_n702), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n806), .A2(new_n807), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n802), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n792), .A2(new_n801), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n789), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n821), .B1(KEYINPUT90), .B2(KEYINPUT36), .C1(new_n824), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n788), .B1(new_n828), .B2(new_n829), .ZN(G311));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n787), .B(KEYINPUT97), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(G150));
  AOI22_X1  g408(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(new_n504), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n512), .A2(G93), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n519), .A2(G55), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n541), .B(new_n542), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT98), .A4(new_n539), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(KEYINPUT98), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n545), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT38), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n631), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n850), .A2(new_n851), .A3(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n838), .A2(G860), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n815), .B(new_n646), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n482), .A2(G142), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n484), .A2(G130), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n469), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n498), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n762), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n752), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n752), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(new_n710), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n868), .A2(new_n752), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n711), .B1(new_n873), .B2(new_n869), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n856), .B(new_n865), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n873), .B(new_n869), .C1(new_n709), .C2(new_n707), .ZN(new_n876));
  INV_X1    g451(.A(new_n711), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n870), .B2(new_n871), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n857), .A2(new_n862), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n857), .A2(new_n862), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n856), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n863), .A2(KEYINPUT101), .A3(new_n864), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n876), .A2(new_n878), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n643), .A2(new_n488), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n643), .A2(new_n488), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(G160), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n889), .B2(new_n890), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n884), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n894), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n875), .A2(new_n899), .A3(new_n883), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n875), .A2(new_n883), .A3(KEYINPUT102), .A4(new_n899), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g480(.A1(new_n838), .A2(G868), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(G288), .ZN(new_n907));
  NOR2_X1   g482(.A1(G305), .A2(new_n603), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G305), .A2(new_n603), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(new_n907), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n912), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n627), .B2(new_n614), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n627), .A2(new_n919), .A3(new_n614), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(G299), .B2(new_n631), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n614), .B(new_n562), .C1(new_n570), .C2(new_n571), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT41), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n919), .B1(new_n627), .B2(new_n614), .ZN(new_n926));
  NAND3_X1  g501(.A1(G299), .A2(KEYINPUT104), .A3(new_n631), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n627), .A2(new_n614), .ZN(new_n931));
  INV_X1    g506(.A(new_n924), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n917), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n635), .B(new_n846), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n924), .B1(new_n920), .B2(new_n921), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n916), .A2(KEYINPUT106), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n911), .A2(new_n914), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n937), .A4(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n906), .B1(new_n947), .B2(G868), .ZN(G295));
  AOI21_X1  g523(.A(new_n906), .B1(new_n947), .B2(G868), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  AOI21_X1  g527(.A(G286), .B1(new_n574), .B2(new_n575), .ZN(new_n953));
  NOR2_X1   g528(.A1(G171), .A2(G168), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n846), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n841), .B(new_n845), .C1(new_n953), .C2(new_n954), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n933), .B1(new_n928), .B2(new_n929), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT105), .B(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n952), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n932), .B1(new_n926), .B2(new_n927), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n957), .B2(new_n956), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n952), .B1(new_n934), .B2(new_n958), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(new_n966), .A3(new_n941), .ZN(new_n967));
  INV_X1    g542(.A(G37), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n938), .A2(KEYINPUT108), .A3(new_n917), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n962), .B2(KEYINPUT41), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n918), .B1(new_n627), .B2(new_n614), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n963), .B1(new_n973), .B2(new_n958), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n974), .B2(new_n915), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n951), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n973), .A2(new_n958), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n941), .B1(new_n977), .B2(new_n963), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(new_n915), .A3(new_n961), .A4(new_n964), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n978), .A2(new_n981), .A3(KEYINPUT109), .A4(new_n968), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n950), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n967), .A2(G37), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n941), .B1(new_n965), .B2(new_n966), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT43), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT44), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n950), .B1(new_n984), .B2(new_n985), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n967), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(G397));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n498), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n482), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n476), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT67), .B1(new_n476), .B2(G2105), .ZN(new_n999));
  OAI211_X1 g574(.A(G40), .B(new_n997), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n762), .B(new_n764), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n752), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1001), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1006), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1005), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n1011), .B(KEYINPUT47), .Z(new_n1012));
  NAND3_X1  g587(.A1(new_n1001), .A2(G1996), .A3(new_n1004), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1003), .B1(new_n1009), .B2(new_n752), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1015), .B(new_n1016), .C1(new_n1006), .C2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n815), .B(new_n818), .Z(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1001), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n603), .A2(new_n1001), .A3(new_n805), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1023));
  OR2_X1    g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n816), .A2(new_n818), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1018), .A2(new_n1027), .B1(G2067), .B2(new_n762), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1012), .B(new_n1026), .C1(new_n1001), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1384), .B1(new_n495), .B2(new_n497), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g606(.A(G160), .B(G40), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT115), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1000), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1033), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n996), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1971), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1041), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1056), .B2(new_n1042), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1055), .B(new_n1052), .C1(new_n1057), .C2(new_n1047), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1036), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1046), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(G8), .A3(new_n1053), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  INV_X1    g638(.A(new_n591), .ZN(new_n1064));
  AOI211_X1 g639(.A(G1981), .B(new_n1064), .C1(new_n587), .C2(new_n589), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n1064), .B2(new_n586), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT49), .B(new_n1066), .C1(G305), .C2(G1981), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n994), .A2(new_n1000), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1049), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT112), .B(G8), .C1(new_n994), .C2(new_n1000), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n797), .A2(G1976), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  INV_X1    g653(.A(G1976), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(G288), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1074), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1062), .A2(new_n1075), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1054), .A2(new_n1058), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1000), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1033), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT125), .B(G1961), .Z(new_n1087));
  INV_X1    g662(.A(G2078), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n996), .A2(new_n1088), .A3(new_n1039), .A4(new_n1043), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1086), .A2(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(G301), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n472), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n996), .A2(new_n477), .A3(new_n1043), .A4(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT54), .B(new_n1093), .C1(new_n1097), .C2(new_n537), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1102));
  AND4_X1   g677(.A1(G301), .A2(new_n1101), .A3(new_n1102), .A4(new_n1096), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G2084), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1037), .A2(new_n1106), .A3(new_n1039), .A4(new_n1033), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1966), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1044), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1085), .A2(KEYINPUT118), .A3(new_n1106), .A4(new_n1033), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .A4(G168), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1113), .A2(new_n1114), .A3(G8), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1112), .A3(new_n1111), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G286), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(G8), .A3(new_n1113), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(KEYINPUT51), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1105), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1044), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1086), .A2(new_n742), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n562), .A2(new_n1126), .A3(new_n565), .A4(new_n569), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n627), .B2(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT120), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1127), .B(new_n1130), .C1(new_n627), .C2(new_n1126), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1125), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n1129), .A3(new_n1124), .A4(new_n1131), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1086), .A2(new_n784), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1071), .A2(new_n764), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n631), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n631), .B2(KEYINPUT124), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1138), .B(new_n1142), .C1(new_n1059), .C2(G1348), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n614), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n614), .A2(new_n1144), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1137), .A2(new_n1138), .A3(new_n1142), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n996), .A2(new_n1009), .A3(new_n1039), .A4(new_n1043), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n994), .B2(new_n1000), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n545), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1153), .B(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(KEYINPUT61), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1149), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(new_n1136), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1135), .B(new_n1140), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1120), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1119), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1113), .A2(G8), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1114), .B1(new_n1166), .B2(new_n1117), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT62), .B1(new_n1167), .B2(new_n1115), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(new_n1100), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1084), .B1(new_n1163), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1059), .A2(new_n1036), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1052), .B1(new_n1171), .B2(new_n1049), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G286), .A2(new_n1049), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(KEYINPUT63), .A3(new_n1116), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1083), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT119), .B1(new_n1082), .B2(new_n1174), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1116), .A2(new_n1173), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1054), .A2(new_n1058), .A3(new_n1083), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1065), .B(KEYINPUT113), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n797), .A2(new_n1079), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT114), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1075), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1074), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1075), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1188), .A2(new_n1189), .B1(new_n1190), .B2(new_n1062), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1170), .A2(new_n1184), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(G290), .A2(G1986), .A3(new_n1001), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1021), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT110), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1020), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1029), .B1(new_n1192), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g772(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1199), .B1(new_n666), .B2(new_n668), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n904), .B(new_n1200), .C1(new_n989), .C2(new_n990), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


