//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G226gat), .A2(G233gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT29), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n220), .B(new_n221), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT64), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT27), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G183gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT28), .A4(new_n224), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT28), .A4(new_n224), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(G190gat), .B1(new_n233), .B2(new_n241), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n237), .B(new_n240), .C1(new_n245), .C2(KEYINPUT28), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n215), .A2(KEYINPUT26), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n214), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n218), .A2(new_n251), .B1(new_n215), .B2(KEYINPUT26), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n250), .A2(new_n252), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n232), .B1(new_n246), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n228), .B(KEYINPUT65), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n230), .B(new_n220), .C1(new_n255), .C2(new_n227), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT25), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n213), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n238), .A2(new_n241), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT28), .B1(new_n259), .B2(new_n243), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n240), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n232), .ZN(new_n263));
  AND4_X1   g062(.A1(new_n210), .A2(new_n262), .A3(new_n257), .A4(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n209), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT75), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n257), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n212), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n254), .A2(new_n210), .A3(new_n257), .ZN(new_n269));
  INV_X1    g068(.A(new_n208), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n207), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n265), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT75), .B(new_n209), .C1(new_n258), .C2(new_n264), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT76), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G8gat), .ZN(new_n278));
  INV_X1    g077(.A(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT30), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G141gat), .B(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(KEYINPUT2), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n292), .C1(new_n288), .C2(KEYINPUT2), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(G127gat), .A2(G134gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(G127gat), .A2(G134gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT69), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  INV_X1    g101(.A(G134gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g104(.A1(G127gat), .A2(G134gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT1), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT70), .B(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n310), .B1(new_n315), .B2(new_n309), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n299), .B2(new_n300), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n304), .A2(new_n318), .A3(new_n306), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT73), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n316), .A2(new_n320), .A3(new_n324), .A4(new_n321), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n298), .B(new_n314), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n314), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT70), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G113gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n330));
  OAI21_X1  g129(.A(G120gat), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n331), .A2(new_n310), .B1(new_n317), .B2(new_n319), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n324), .B1(new_n332), .B2(new_n321), .ZN(new_n333));
  AND4_X1   g132(.A1(new_n324), .A2(new_n316), .A3(new_n320), .A4(new_n321), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n327), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n298), .B(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n326), .A2(KEYINPUT4), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n314), .B1(new_n323), .B2(new_n325), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n298), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n338), .B(new_n341), .C1(new_n346), .C2(KEYINPUT4), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT0), .B(G57gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g150(.A(new_n298), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n298), .B(KEYINPUT3), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT4), .B(new_n339), .C1(new_n354), .C2(new_n343), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n346), .A2(KEYINPUT4), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n343), .A2(new_n352), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n340), .B1(new_n357), .B2(new_n326), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n347), .B(new_n351), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n353), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n343), .A2(new_n344), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT74), .B(new_n314), .C1(new_n323), .C2(new_n325), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n352), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n335), .A2(new_n298), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n353), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n371), .B2(new_n340), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n351), .B1(new_n373), .B2(new_n347), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n362), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n347), .B1(new_n356), .B2(new_n359), .ZN(new_n376));
  INV_X1    g175(.A(new_n351), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n287), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n267), .B1(new_n364), .B2(new_n365), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n262), .A2(new_n257), .A3(new_n263), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n342), .A3(new_n345), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n382), .A2(new_n384), .A3(G227gat), .A4(G233gat), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n385), .A2(KEYINPUT32), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n384), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT34), .ZN(new_n388));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n387), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT34), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n385), .A2(KEYINPUT32), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G15gat), .B(G43gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  AND2_X1   g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n392), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n209), .A2(KEYINPUT29), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n271), .A2(new_n211), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT77), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n352), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n211), .B1(new_n298), .B2(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n209), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n412), .A2(new_n209), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n352), .B1(new_n409), .B2(new_n336), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI22_X1  g217(.A1(new_n411), .A2(new_n415), .B1(new_n418), .B2(new_n414), .ZN(new_n419));
  XOR2_X1   g218(.A(G78gat), .B(G106gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT31), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n421), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n403), .B1(new_n392), .B2(new_n397), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n405), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT35), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(KEYINPUT83), .A2(KEYINPUT35), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n381), .A2(new_n429), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n425), .A2(new_n426), .ZN(new_n435));
  INV_X1    g234(.A(new_n403), .ZN(new_n436));
  INV_X1    g235(.A(new_n397), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n396), .B1(new_n394), .B2(new_n395), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n439), .A3(new_n404), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n284), .A2(new_n286), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n379), .B2(new_n375), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n430), .B(new_n431), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n275), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n265), .A2(KEYINPUT81), .A3(new_n272), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(KEYINPUT37), .C1(KEYINPUT81), .C2(new_n265), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .A4(new_n280), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n380), .A2(KEYINPUT82), .A3(new_n282), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n446), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n280), .B1(new_n275), .B2(new_n445), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT38), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n376), .A2(new_n377), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n361), .A3(new_n360), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n450), .A2(new_n456), .A3(new_n378), .A4(new_n282), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n370), .A2(new_n353), .A3(new_n339), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n353), .A2(new_n367), .B1(new_n343), .B2(new_n354), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n366), .B2(new_n367), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT39), .B(new_n461), .C1(new_n463), .C2(new_n339), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n338), .B1(new_n346), .B2(KEYINPUT4), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n340), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n464), .A2(new_n467), .A3(KEYINPUT40), .A4(new_n351), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n284), .A2(new_n468), .A3(new_n455), .A4(new_n286), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n464), .A2(new_n351), .A3(new_n467), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT79), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n472), .A2(KEYINPUT79), .A3(new_n473), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n470), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT80), .B1(new_n477), .B2(new_n469), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n460), .A2(new_n435), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n405), .A2(new_n428), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n405), .B2(new_n428), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n427), .B(KEYINPUT78), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n481), .A2(new_n483), .B1(new_n484), .B2(new_n442), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n444), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G127gat), .B(G155gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(new_n204), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(G1gat), .ZN(new_n491));
  INV_X1    g290(.A(G1gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(KEYINPUT87), .A3(KEYINPUT16), .ZN(new_n493));
  OR2_X1    g292(.A1(G15gat), .A2(G22gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(G15gat), .A2(G22gat), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n491), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n492), .A3(new_n495), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n492), .A2(KEYINPUT87), .A3(KEYINPUT16), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT87), .B1(new_n492), .B2(KEYINPUT16), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n498), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G8gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT89), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n496), .B2(new_n498), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n494), .A2(new_n492), .A3(new_n495), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT88), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n506), .A3(new_n509), .ZN(new_n514));
  NAND2_X1  g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT9), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(G57gat), .A2(G64gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(G57gat), .A2(G64gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(KEYINPUT92), .A3(new_n516), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n519), .A2(new_n522), .A3(new_n525), .A4(new_n523), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(G183gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(G183gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n532), .B2(new_n533), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n488), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  INV_X1    g339(.A(new_n488), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n544), .B(new_n545), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n539), .A2(new_n542), .A3(new_n546), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G50gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT86), .B1(new_n552), .B2(G43gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556));
  INV_X1    g355(.A(G29gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n279), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n279), .A2(KEYINPUT85), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n563), .A3(G29gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n555), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT85), .B(G36gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n567), .A2(G29gat), .B1(new_n558), .B2(new_n559), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n565), .B(new_n566), .C1(new_n568), .C2(KEYINPUT15), .ZN(new_n569));
  INV_X1    g368(.A(new_n566), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n570), .A3(new_n555), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n576), .A2(new_n579), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n569), .A2(KEYINPUT17), .A3(new_n571), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n574), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT93), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT41), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n584), .B(new_n585), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n572), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n224), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n224), .B1(new_n589), .B2(new_n595), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n205), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(G218gat), .A3(new_n596), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n591), .A2(new_n592), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n291), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT94), .B(G134gat), .Z(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n603), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n551), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n486), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n574), .A2(new_n513), .A3(new_n514), .A4(new_n588), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n511), .B1(new_n507), .B2(new_n510), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n514), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n572), .ZN(new_n618));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT18), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n614), .A2(new_n618), .A3(new_n622), .A4(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT90), .ZN(new_n625));
  INV_X1    g424(.A(new_n572), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n513), .A2(new_n626), .A3(new_n514), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n618), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n619), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n617), .A2(KEYINPUT90), .A3(new_n572), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G113gat), .B(G141gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G169gat), .B(G197gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n613), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n628), .A2(new_n631), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n642), .A2(new_n630), .B1(new_n621), .B2(new_n623), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(KEYINPUT91), .A3(new_n639), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n641), .A2(new_n644), .B1(new_n633), .B2(new_n640), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n217), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(G204gat), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n584), .A2(KEYINPUT96), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n594), .A2(new_n527), .A3(new_n528), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n527), .A2(new_n528), .A3(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n587), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n649), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n650), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n652), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n529), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI211_X1 g461(.A(KEYINPUT97), .B(new_n650), .C1(new_n652), .C2(new_n654), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n657), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n648), .B1(new_n662), .B2(new_n655), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT98), .B(new_n648), .C1(new_n662), .C2(new_n655), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT99), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n645), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n612), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n380), .A2(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n380), .A2(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n492), .ZN(G1324gat));
  NOR2_X1   g477(.A1(new_n672), .A2(new_n441), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n490), .A2(new_n506), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n490), .A2(new_n506), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n679), .A2(KEYINPUT42), .A3(new_n681), .A4(new_n682), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n685), .B(new_n686), .C1(new_n506), .C2(new_n679), .ZN(G1325gat));
  INV_X1    g486(.A(new_n672), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n481), .A2(new_n483), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT101), .Z(new_n690));
  AND3_X1   g489(.A1(new_n688), .A2(G15gat), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(G15gat), .B1(new_n688), .B2(new_n480), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1326gat));
  INV_X1    g492(.A(new_n484), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n672), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT102), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n695), .B(new_n697), .ZN(G1327gat));
  NAND2_X1  g497(.A1(new_n479), .A2(new_n485), .ZN(new_n699));
  INV_X1    g498(.A(new_n444), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(KEYINPUT44), .A3(new_n609), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n603), .B(new_n607), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n486), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n667), .A2(new_n668), .ZN(new_n706));
  INV_X1    g505(.A(new_n664), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT99), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT99), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n709), .B(new_n664), .C1(new_n667), .C2(new_n668), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT104), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n550), .A2(new_n645), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n702), .A2(new_n705), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n715), .A2(new_n716), .A3(new_n676), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n715), .B2(new_n676), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(G29gat), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n711), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n486), .A2(new_n704), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n557), .A3(new_n675), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n724), .ZN(G1328gat));
  NOR2_X1   g524(.A1(new_n441), .A2(new_n567), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n567), .B1(new_n715), .B2(new_n441), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(KEYINPUT106), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(G1329gat));
  OAI21_X1  g532(.A(G43gat), .B1(new_n715), .B2(new_n689), .ZN(new_n734));
  INV_X1    g533(.A(new_n480), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(KEYINPUT47), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n701), .B2(new_n609), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n486), .A2(new_n703), .A3(new_n704), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n742), .A2(new_n690), .A3(new_n713), .A4(new_n714), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n743), .B2(G43gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n738), .B1(new_n744), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n486), .A2(new_n704), .ZN(new_n747));
  INV_X1    g546(.A(new_n720), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n484), .A2(new_n552), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n486), .A2(KEYINPUT107), .A3(new_n704), .A4(new_n720), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G50gat), .B1(new_n715), .B2(new_n435), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT48), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n742), .A2(new_n484), .A3(new_n713), .A4(new_n714), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g557(.A1(new_n633), .A2(new_n640), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT91), .B1(new_n643), .B2(new_n639), .ZN(new_n760));
  AND4_X1   g559(.A1(KEYINPUT91), .A2(new_n624), .A3(new_n632), .A4(new_n639), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n486), .A2(new_n762), .A3(new_n611), .A4(new_n713), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n675), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NAND4_X1  g564(.A1(new_n701), .A2(new_n645), .A3(new_n610), .A4(new_n712), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n441), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n763), .A2(G71gat), .A3(new_n690), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n766), .A2(new_n735), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(G71gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n763), .A2(new_n484), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n550), .A2(new_n762), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n747), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  INV_X1    g579(.A(new_n778), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n486), .A2(new_n780), .A3(new_n704), .A4(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(new_n580), .A3(new_n675), .A4(new_n670), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n781), .A2(new_n711), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n742), .A2(new_n675), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n580), .B2(new_n786), .ZN(G1336gat));
  NAND3_X1  g586(.A1(new_n712), .A2(new_n581), .A3(new_n287), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT108), .Z(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n779), .B2(new_n782), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n702), .A2(new_n705), .A3(new_n287), .A4(new_n785), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n789), .B(KEYINPUT109), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n783), .A2(new_n795), .B1(G92gat), .B2(new_n791), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n793), .ZN(G1337gat));
  NOR2_X1   g596(.A1(new_n735), .A2(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n670), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n742), .A2(new_n690), .A3(new_n785), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G99gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1338gat));
  NOR2_X1   g601(.A1(new_n713), .A2(G106gat), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n427), .B(new_n803), .C1(new_n779), .C2(new_n782), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n702), .A2(new_n705), .A3(new_n484), .A4(new_n785), .ZN(new_n805));
  XNOR2_X1  g604(.A(KEYINPUT110), .B(G106gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n702), .A2(new_n705), .A3(new_n427), .A4(new_n785), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n806), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n804), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(G1339gat));
  NAND4_X1  g613(.A1(new_n550), .A2(new_n645), .A3(new_n711), .A4(new_n704), .ZN(new_n815));
  INV_X1    g614(.A(new_n638), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n614), .A2(new_n618), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n642), .A2(new_n630), .B1(new_n619), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n641), .A2(new_n644), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n609), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n660), .A2(new_n658), .A3(new_n661), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n821), .A2(new_n662), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n662), .A2(new_n822), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT112), .B1(new_n824), .B2(new_n648), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n826), .B(new_n649), .C1(new_n662), .C2(new_n822), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(KEYINPUT55), .B(new_n823), .C1(new_n825), .C2(new_n827), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT113), .A3(new_n707), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT113), .B1(new_n831), .B2(new_n707), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n820), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n762), .B(new_n830), .C1(new_n833), .C2(new_n832), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n816), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n760), .B2(new_n761), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n839), .B2(new_n711), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n819), .A2(new_n670), .A3(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n835), .B1(new_n842), .B2(new_n704), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n815), .B1(new_n843), .B2(new_n550), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n676), .A2(new_n287), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n429), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n762), .C1(new_n329), .C2(new_n330), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n844), .A2(new_n850), .A3(new_n694), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n844), .B2(new_n694), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n735), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n762), .A3(new_n845), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n854), .B2(G113gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n844), .A2(new_n694), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT115), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n844), .A2(new_n850), .A3(new_n694), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n857), .A2(new_n480), .A3(new_n845), .A4(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n849), .B(G113gat), .C1(new_n859), .C2(new_n645), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n848), .B1(new_n855), .B2(new_n861), .ZN(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n859), .B2(new_n713), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n309), .A3(new_n670), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1341gat));
  NAND4_X1  g664(.A1(new_n853), .A2(G127gat), .A3(new_n550), .A4(new_n845), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n859), .A2(new_n302), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n550), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n847), .A2(new_n550), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n302), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n867), .A2(new_n870), .A3(new_n872), .ZN(G1342gat));
  NAND3_X1  g672(.A1(new_n847), .A2(new_n303), .A3(new_n609), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n859), .B2(new_n704), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n690), .A2(new_n435), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n846), .ZN(new_n880));
  INV_X1    g679(.A(G141gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n762), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n839), .B2(new_n711), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n819), .A2(new_n670), .A3(KEYINPUT118), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n831), .A2(new_n707), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n762), .A2(new_n830), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n835), .B1(new_n888), .B2(new_n704), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n815), .B1(new_n889), .B2(new_n550), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n484), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n845), .A2(new_n689), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n844), .A2(new_n894), .A3(new_n427), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n645), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1344gat));
  NAND4_X1  g701(.A1(new_n892), .A2(new_n670), .A3(new_n893), .A4(new_n895), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(KEYINPUT59), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n903), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n844), .A2(new_n427), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT57), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n815), .B(KEYINPUT121), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n889), .B2(new_n550), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n894), .A3(new_n484), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n910), .A2(new_n670), .A3(new_n893), .A4(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(G148gat), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n907), .A2(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n880), .A2(new_n905), .A3(new_n670), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1345gat));
  NOR3_X1   g718(.A1(new_n896), .A2(new_n290), .A3(new_n551), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n879), .A2(new_n846), .A3(new_n550), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT122), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n290), .ZN(G1346gat));
  AND4_X1   g722(.A1(new_n291), .A2(new_n879), .A3(new_n846), .A4(new_n609), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT123), .ZN(new_n925));
  OAI21_X1  g724(.A(G162gat), .B1(new_n896), .B2(new_n704), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  AND2_X1   g726(.A1(new_n844), .A2(new_n676), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n440), .A2(new_n441), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n216), .A3(new_n762), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n676), .A2(new_n287), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT124), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n853), .A2(new_n762), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n935), .B2(G169gat), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n857), .A2(new_n480), .A3(new_n858), .A4(new_n934), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(G169gat), .C1(new_n937), .C2(new_n645), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n931), .B1(new_n936), .B2(new_n939), .ZN(G1348gat));
  NOR3_X1   g739(.A1(new_n937), .A2(new_n217), .A3(new_n713), .ZN(new_n941));
  AOI21_X1  g740(.A(G176gat), .B1(new_n930), .B2(new_n670), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n937), .B2(new_n551), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n550), .A3(new_n238), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT60), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1350gat));
  NAND4_X1  g749(.A1(new_n928), .A2(new_n224), .A3(new_n609), .A4(new_n929), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT126), .Z(new_n952));
  OAI21_X1  g751(.A(G190gat), .B1(new_n937), .B2(new_n704), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g754(.A(KEYINPUT61), .B(G190gat), .C1(new_n937), .C2(new_n704), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(G1351gat));
  INV_X1    g756(.A(new_n690), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n910), .A2(new_n958), .A3(new_n913), .A4(new_n934), .ZN(new_n959));
  OAI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n645), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n879), .A2(new_n928), .A3(new_n287), .ZN(new_n961));
  INV_X1    g760(.A(G197gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n962), .A3(new_n762), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(G1352gat));
  XOR2_X1   g763(.A(KEYINPUT127), .B(G204gat), .Z(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n961), .A2(new_n670), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n959), .B2(new_n713), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n961), .A2(new_n970), .A3(new_n670), .A4(new_n966), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n961), .A2(new_n204), .A3(new_n550), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n912), .A2(new_n894), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n974), .A2(new_n484), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n975), .A2(new_n550), .A3(new_n958), .A4(new_n934), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n977));
  OAI211_X1 g776(.A(KEYINPUT63), .B(G211gat), .C1(new_n959), .C2(new_n551), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n959), .B2(new_n704), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n205), .A3(new_n609), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


