

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744;

  BUF_X1 U367 ( .A(n708), .Z(n348) );
  AND2_X1 U368 ( .A1(n443), .A2(n440), .ZN(n439) );
  XNOR2_X1 U369 ( .A(n475), .B(n421), .ZN(n677) );
  NOR2_X1 U370 ( .A1(G902), .A2(n625), .ZN(n475) );
  XNOR2_X1 U371 ( .A(n455), .B(G128), .ZN(n505) );
  NAND2_X1 U372 ( .A1(n542), .A2(n361), .ZN(n448) );
  XNOR2_X1 U373 ( .A(n539), .B(n364), .ZN(n542) );
  XNOR2_X1 U374 ( .A(n519), .B(KEYINPUT31), .ZN(n650) );
  NOR2_X1 U375 ( .A1(G902), .A2(n699), .ZN(n501) );
  XNOR2_X2 U376 ( .A(G110), .B(G104), .ZN(n382) );
  XNOR2_X2 U377 ( .A(n433), .B(n554), .ZN(n558) );
  INV_X1 U378 ( .A(n571), .ZN(n347) );
  XOR2_X1 U379 ( .A(n559), .B(KEYINPUT6), .Z(n571) );
  INV_X1 U380 ( .A(KEYINPUT77), .ZN(n384) );
  INV_X1 U381 ( .A(KEYINPUT74), .ZN(n352) );
  INV_X1 U382 ( .A(G143), .ZN(n455) );
  AND2_X1 U383 ( .A1(n412), .A2(n429), .ZN(n408) );
  BUF_X1 U384 ( .A(n550), .Z(n540) );
  XNOR2_X1 U385 ( .A(n397), .B(n518), .ZN(n550) );
  NOR2_X1 U386 ( .A1(n559), .A2(n537), .ZN(n502) );
  NAND2_X1 U387 ( .A1(n597), .A2(n516), .ZN(n397) );
  XNOR2_X1 U388 ( .A(n493), .B(n415), .ZN(n572) );
  XNOR2_X1 U389 ( .A(n505), .B(n467), .ZN(n528) );
  XNOR2_X1 U390 ( .A(n553), .B(KEYINPUT75), .ZN(n554) );
  INV_X1 U391 ( .A(n559), .ZN(n349) );
  AND2_X1 U392 ( .A1(n379), .A2(n730), .ZN(n658) );
  BUF_X1 U393 ( .A(n396), .Z(n350) );
  NAND2_X1 U394 ( .A1(n716), .A2(KEYINPUT74), .ZN(n353) );
  NAND2_X1 U395 ( .A1(n351), .A2(n352), .ZN(n354) );
  NAND2_X1 U396 ( .A1(n353), .A2(n354), .ZN(n506) );
  INV_X1 U397 ( .A(n716), .ZN(n351) );
  XNOR2_X2 U398 ( .A(n569), .B(KEYINPUT45), .ZN(n379) );
  XNOR2_X1 U399 ( .A(n557), .B(n556), .ZN(n396) );
  XNOR2_X1 U400 ( .A(n374), .B(n494), .ZN(n716) );
  NAND2_X1 U401 ( .A1(n406), .A2(n405), .ZN(n557) );
  XNOR2_X1 U402 ( .A(n382), .B(n384), .ZN(n374) );
  NAND2_X1 U403 ( .A1(n432), .A2(n431), .ZN(n433) );
  INV_X1 U404 ( .A(n546), .ZN(n442) );
  XNOR2_X1 U405 ( .A(G902), .B(KEYINPUT15), .ZN(n570) );
  XNOR2_X1 U406 ( .A(n545), .B(KEYINPUT35), .ZN(n546) );
  XNOR2_X1 U407 ( .A(n728), .B(G146), .ZN(n499) );
  XOR2_X1 U408 ( .A(G146), .B(G125), .Z(n503) );
  NOR2_X1 U409 ( .A1(n551), .A2(n572), .ZN(n671) );
  XNOR2_X1 U410 ( .A(n503), .B(n385), .ZN(n726) );
  INV_X1 U411 ( .A(KEYINPUT10), .ZN(n385) );
  NOR2_X1 U412 ( .A1(G953), .A2(G237), .ZN(n468) );
  XOR2_X1 U413 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n460) );
  INV_X1 U414 ( .A(G224), .ZN(n377) );
  AND2_X1 U415 ( .A1(n446), .A2(n599), .ZN(n445) );
  NAND2_X1 U416 ( .A1(n540), .A2(n447), .ZN(n446) );
  XNOR2_X1 U417 ( .A(n485), .B(n486), .ZN(n523) );
  XNOR2_X1 U418 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n485) );
  AND2_X1 U419 ( .A1(n730), .A2(n367), .ZN(n401) );
  NAND2_X1 U420 ( .A1(n549), .A2(n548), .ZN(n664) );
  NOR2_X1 U421 ( .A1(n543), .A2(n442), .ZN(n441) );
  AND2_X1 U422 ( .A1(n437), .A2(n442), .ZN(n436) );
  NAND2_X1 U423 ( .A1(n582), .A2(n661), .ZN(n383) );
  XNOR2_X1 U424 ( .A(n473), .B(n508), .ZN(n474) );
  XNOR2_X1 U425 ( .A(n423), .B(n422), .ZN(n473) );
  XNOR2_X1 U426 ( .A(n470), .B(G101), .ZN(n422) );
  BUF_X1 U427 ( .A(n520), .Z(n591) );
  XNOR2_X1 U428 ( .A(G128), .B(G119), .ZN(n479) );
  XNOR2_X1 U429 ( .A(n414), .B(n484), .ZN(n488) );
  XNOR2_X1 U430 ( .A(n483), .B(n356), .ZN(n414) );
  INV_X1 U431 ( .A(G134), .ZN(n467) );
  NAND2_X1 U432 ( .A1(n523), .A2(G217), .ZN(n395) );
  XNOR2_X1 U433 ( .A(n524), .B(n394), .ZN(n393) );
  INV_X1 U434 ( .A(KEYINPUT9), .ZN(n394) );
  XNOR2_X1 U435 ( .A(n463), .B(n359), .ZN(n411) );
  XNOR2_X1 U436 ( .A(n589), .B(KEYINPUT39), .ZN(n610) );
  BUF_X1 U437 ( .A(n670), .Z(n409) );
  INV_X1 U438 ( .A(n677), .ZN(n559) );
  XNOR2_X1 U439 ( .A(n492), .B(n357), .ZN(n415) );
  INV_X1 U440 ( .A(KEYINPUT47), .ZN(n386) );
  INV_X1 U441 ( .A(KEYINPUT65), .ZN(n430) );
  AND2_X1 U442 ( .A1(n547), .A2(n741), .ZN(n429) );
  XNOR2_X1 U443 ( .A(n509), .B(n456), .ZN(n582) );
  XNOR2_X1 U444 ( .A(n469), .B(n424), .ZN(n423) );
  AND2_X1 U445 ( .A1(n468), .A2(G210), .ZN(n424) );
  XNOR2_X1 U446 ( .A(n501), .B(n500), .ZN(n520) );
  AND2_X1 U447 ( .A1(n552), .A2(n434), .ZN(n431) );
  INV_X1 U448 ( .A(n551), .ZN(n434) );
  XNOR2_X1 U449 ( .A(n454), .B(n528), .ZN(n728) );
  XNOR2_X1 U450 ( .A(n504), .B(G137), .ZN(n454) );
  XNOR2_X1 U451 ( .A(G143), .B(G113), .ZN(n457) );
  XNOR2_X1 U452 ( .A(n388), .B(n459), .ZN(n463) );
  XNOR2_X1 U453 ( .A(n460), .B(n389), .ZN(n388) );
  INV_X1 U454 ( .A(KEYINPUT102), .ZN(n389) );
  XNOR2_X1 U455 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n504) );
  XNOR2_X1 U456 ( .A(n376), .B(n378), .ZN(n373) );
  NOR2_X1 U457 ( .A1(n377), .A2(G953), .ZN(n376) );
  XNOR2_X1 U458 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n378) );
  NOR2_X1 U459 ( .A1(n674), .A2(n578), .ZN(n579) );
  XNOR2_X1 U460 ( .A(n520), .B(KEYINPUT1), .ZN(n670) );
  XNOR2_X1 U461 ( .A(n517), .B(KEYINPUT0), .ZN(n518) );
  AND2_X1 U462 ( .A1(n416), .A2(n362), .ZN(n730) );
  XNOR2_X1 U463 ( .A(G116), .B(G113), .ZN(n471) );
  NAND2_X1 U464 ( .A1(n658), .A2(KEYINPUT2), .ZN(n622) );
  XNOR2_X1 U465 ( .A(n375), .B(n715), .ZN(n698) );
  XNOR2_X1 U466 ( .A(n506), .B(n370), .ZN(n375) );
  XNOR2_X1 U467 ( .A(n372), .B(n371), .ZN(n370) );
  XNOR2_X1 U468 ( .A(n503), .B(n504), .ZN(n371) );
  OR2_X1 U469 ( .A1(n392), .A2(n648), .ZN(n605) );
  NAND2_X1 U470 ( .A1(n347), .A2(n592), .ZN(n392) );
  NAND2_X1 U471 ( .A1(n439), .A2(n435), .ZN(n742) );
  NAND2_X1 U472 ( .A1(n438), .A2(n436), .ZN(n435) );
  NOR2_X1 U473 ( .A1(n587), .A2(n586), .ZN(n600) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n585) );
  INV_X1 U475 ( .A(KEYINPUT30), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n533), .B(n358), .ZN(n549) );
  NOR2_X1 U477 ( .A1(n534), .A2(n549), .ZN(n611) );
  INV_X1 U478 ( .A(G472), .ZN(n421) );
  INV_X1 U479 ( .A(G953), .ZN(n731) );
  XNOR2_X1 U480 ( .A(n726), .B(n480), .ZN(n490) );
  XNOR2_X1 U481 ( .A(G116), .B(G107), .ZN(n525) );
  XNOR2_X1 U482 ( .A(n395), .B(n393), .ZN(n526) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n740) );
  XNOR2_X1 U484 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n417) );
  NAND2_X1 U485 ( .A1(n610), .A2(n611), .ZN(n418) );
  BUF_X1 U486 ( .A(n742), .Z(n407) );
  XNOR2_X1 U487 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n556) );
  XNOR2_X1 U488 ( .A(n611), .B(KEYINPUT109), .ZN(n648) );
  INV_X1 U489 ( .A(KEYINPUT56), .ZN(n449) );
  XOR2_X1 U490 ( .A(n381), .B(n368), .Z(n355) );
  XOR2_X1 U491 ( .A(G140), .B(KEYINPUT84), .Z(n356) );
  XOR2_X1 U492 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n357) );
  XOR2_X1 U493 ( .A(n531), .B(n530), .Z(n358) );
  XOR2_X1 U494 ( .A(n458), .B(n457), .Z(n359) );
  XOR2_X1 U495 ( .A(G119), .B(KEYINPUT3), .Z(n360) );
  AND2_X1 U496 ( .A1(n541), .A2(n543), .ZN(n361) );
  AND2_X1 U497 ( .A1(n657), .A2(n656), .ZN(n362) );
  NAND2_X1 U498 ( .A1(n572), .A2(n409), .ZN(n363) );
  XNOR2_X1 U499 ( .A(KEYINPUT92), .B(KEYINPUT33), .ZN(n364) );
  INV_X1 U500 ( .A(n543), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n532), .B(n466), .ZN(n365) );
  NAND2_X1 U502 ( .A1(n619), .A2(KEYINPUT85), .ZN(n403) );
  XOR2_X1 U503 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n366) );
  OR2_X1 U504 ( .A1(n619), .A2(KEYINPUT85), .ZN(n367) );
  INV_X1 U505 ( .A(n714), .ZN(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n368) );
  XOR2_X1 U507 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n369) );
  XNOR2_X1 U508 ( .A(n505), .B(n373), .ZN(n372) );
  NAND2_X1 U509 ( .A1(n698), .A2(n570), .ZN(n509) );
  BUF_X1 U510 ( .A(n716), .Z(n380) );
  BUF_X1 U511 ( .A(G104), .Z(n634) );
  NAND2_X1 U512 ( .A1(n349), .A2(n661), .ZN(n420) );
  BUF_X1 U513 ( .A(n698), .Z(n381) );
  XNOR2_X2 U514 ( .A(n383), .B(KEYINPUT19), .ZN(n597) );
  NOR2_X1 U515 ( .A1(n605), .A2(n383), .ZN(n607) );
  AND2_X2 U516 ( .A1(n624), .A2(n622), .ZN(n708) );
  XNOR2_X1 U517 ( .A(n618), .B(n366), .ZN(n416) );
  NAND2_X1 U518 ( .A1(n654), .A2(n609), .ZN(n391) );
  XNOR2_X1 U519 ( .A(n387), .B(n386), .ZN(n604) );
  NOR2_X1 U520 ( .A1(n646), .A2(n666), .ZN(n387) );
  NAND2_X1 U521 ( .A1(n404), .A2(n621), .ZN(n624) );
  NAND2_X1 U522 ( .A1(n400), .A2(KEYINPUT85), .ZN(n399) );
  XNOR2_X1 U523 ( .A(n462), .B(n411), .ZN(n532) );
  NAND2_X1 U524 ( .A1(n390), .A2(n617), .ZN(n618) );
  XNOR2_X1 U525 ( .A(n391), .B(KEYINPUT71), .ZN(n390) );
  NAND2_X1 U526 ( .A1(n608), .A2(n409), .ZN(n654) );
  NAND2_X1 U527 ( .A1(n396), .A2(n641), .ZN(n565) );
  XNOR2_X1 U528 ( .A(n350), .B(n744), .ZN(G21) );
  NAND2_X1 U529 ( .A1(n398), .A2(n399), .ZN(n402) );
  NAND2_X1 U530 ( .A1(n379), .A2(n403), .ZN(n398) );
  INV_X1 U531 ( .A(n379), .ZN(n400) );
  NAND2_X1 U532 ( .A1(n402), .A2(n401), .ZN(n404) );
  NAND2_X1 U533 ( .A1(n708), .A2(G475), .ZN(n427) );
  NAND2_X1 U534 ( .A1(n708), .A2(G210), .ZN(n453) );
  NOR2_X1 U535 ( .A1(n555), .A2(n363), .ZN(n405) );
  XNOR2_X1 U536 ( .A(n453), .B(n355), .ZN(n452) );
  XNOR2_X1 U537 ( .A(n427), .B(n365), .ZN(n426) );
  INV_X1 U538 ( .A(n558), .ZN(n406) );
  NAND2_X1 U539 ( .A1(n426), .A2(n451), .ZN(n425) );
  NAND2_X1 U540 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U541 ( .A(n425), .B(n369), .ZN(G60) );
  XNOR2_X1 U542 ( .A(n450), .B(n449), .ZN(G51) );
  INV_X1 U543 ( .A(n542), .ZN(n660) );
  NAND2_X1 U544 ( .A1(n410), .A2(n408), .ZN(n428) );
  XNOR2_X1 U545 ( .A(n499), .B(n498), .ZN(n699) );
  XNOR2_X1 U546 ( .A(n561), .B(n430), .ZN(n410) );
  NAND2_X1 U547 ( .A1(n413), .A2(KEYINPUT44), .ZN(n412) );
  INV_X1 U548 ( .A(n742), .ZN(n413) );
  XNOR2_X1 U549 ( .A(n428), .B(KEYINPUT89), .ZN(n568) );
  INV_X1 U550 ( .A(n550), .ZN(n432) );
  NAND2_X1 U551 ( .A1(n660), .A2(n447), .ZN(n437) );
  INV_X1 U552 ( .A(n444), .ZN(n438) );
  NAND2_X1 U553 ( .A1(n660), .A2(n441), .ZN(n440) );
  NAND2_X1 U554 ( .A1(n444), .A2(n546), .ZN(n443) );
  NAND2_X1 U555 ( .A1(n448), .A2(n445), .ZN(n444) );
  NOR2_X1 U556 ( .A1(G952), .A2(n731), .ZN(n714) );
  XNOR2_X1 U557 ( .A(n499), .B(n474), .ZN(n625) );
  AND2_X1 U558 ( .A1(n510), .A2(G210), .ZN(n456) );
  INV_X1 U559 ( .A(KEYINPUT98), .ZN(n478) );
  XNOR2_X1 U560 ( .A(n727), .B(n496), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U562 ( .A(n506), .B(n497), .ZN(n498) );
  INV_X1 U563 ( .A(KEYINPUT62), .ZN(n626) );
  INV_X1 U564 ( .A(G469), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n627), .B(n626), .ZN(n628) );
  INV_X1 U566 ( .A(KEYINPUT123), .ZN(n709) );
  INV_X1 U567 ( .A(KEYINPUT80), .ZN(n545) );
  XNOR2_X1 U568 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U569 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U570 ( .A(n631), .B(KEYINPUT114), .ZN(n632) );
  XNOR2_X1 U571 ( .A(n712), .B(n711), .ZN(n713) );
  XOR2_X1 U572 ( .A(G122), .B(n634), .Z(n458) );
  NAND2_X1 U573 ( .A1(G214), .A2(n468), .ZN(n459) );
  XOR2_X1 U574 ( .A(G131), .B(G140), .Z(n495) );
  INV_X1 U575 ( .A(n495), .ZN(n461) );
  XOR2_X1 U576 ( .A(n461), .B(n726), .Z(n462) );
  XOR2_X1 U577 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n465) );
  XNOR2_X1 U578 ( .A(KEYINPUT94), .B(KEYINPUT68), .ZN(n464) );
  XNOR2_X1 U579 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U580 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n469) );
  XNOR2_X1 U581 ( .A(G131), .B(KEYINPUT100), .ZN(n470) );
  XNOR2_X1 U582 ( .A(n360), .B(n471), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n472), .B(KEYINPUT73), .ZN(n508) );
  NAND2_X1 U584 ( .A1(G234), .A2(n570), .ZN(n476) );
  XNOR2_X1 U585 ( .A(KEYINPUT20), .B(n476), .ZN(n491) );
  NAND2_X1 U586 ( .A1(n491), .A2(G221), .ZN(n477) );
  XOR2_X1 U587 ( .A(KEYINPUT21), .B(n477), .Z(n673) );
  XNOR2_X1 U588 ( .A(KEYINPUT99), .B(n673), .ZN(n551) );
  XOR2_X1 U589 ( .A(KEYINPUT79), .B(KEYINPUT23), .Z(n482) );
  XNOR2_X1 U590 ( .A(G137), .B(G110), .ZN(n481) );
  XNOR2_X1 U591 ( .A(n482), .B(n481), .ZN(n484) );
  XOR2_X1 U592 ( .A(KEYINPUT97), .B(KEYINPUT24), .Z(n483) );
  NAND2_X1 U593 ( .A1(n731), .A2(G234), .ZN(n486) );
  NAND2_X1 U594 ( .A1(G221), .A2(n523), .ZN(n487) );
  XNOR2_X1 U595 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n490), .B(n489), .ZN(n710) );
  NOR2_X1 U597 ( .A1(G902), .A2(n710), .ZN(n493) );
  NAND2_X1 U598 ( .A1(G217), .A2(n491), .ZN(n492) );
  XNOR2_X1 U599 ( .A(G101), .B(G107), .ZN(n494) );
  XOR2_X1 U600 ( .A(KEYINPUT96), .B(n495), .Z(n727) );
  AND2_X1 U601 ( .A1(G227), .A2(n731), .ZN(n496) );
  NAND2_X1 U602 ( .A1(n671), .A2(n670), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT101), .B(n502), .ZN(n682) );
  XNOR2_X1 U604 ( .A(KEYINPUT16), .B(G122), .ZN(n507) );
  XNOR2_X1 U605 ( .A(n508), .B(n507), .ZN(n715) );
  OR2_X1 U606 ( .A1(G237), .A2(G902), .ZN(n510) );
  NAND2_X1 U607 ( .A1(G214), .A2(n510), .ZN(n661) );
  NAND2_X1 U608 ( .A1(G234), .A2(G237), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n511), .B(KEYINPUT14), .ZN(n513) );
  NAND2_X1 U610 ( .A1(G952), .A2(n513), .ZN(n690) );
  NOR2_X1 U611 ( .A1(n690), .A2(G953), .ZN(n512) );
  XNOR2_X1 U612 ( .A(n512), .B(KEYINPUT95), .ZN(n576) );
  NAND2_X1 U613 ( .A1(G902), .A2(n513), .ZN(n573) );
  INV_X1 U614 ( .A(n573), .ZN(n514) );
  NOR2_X1 U615 ( .A1(G898), .A2(n731), .ZN(n717) );
  NAND2_X1 U616 ( .A1(n514), .A2(n717), .ZN(n515) );
  NAND2_X1 U617 ( .A1(n576), .A2(n515), .ZN(n516) );
  INV_X1 U618 ( .A(KEYINPUT91), .ZN(n517) );
  NOR2_X1 U619 ( .A1(n682), .A2(n540), .ZN(n519) );
  NAND2_X1 U620 ( .A1(n591), .A2(n671), .ZN(n587) );
  INV_X1 U621 ( .A(n587), .ZN(n522) );
  NOR2_X1 U622 ( .A1(n349), .A2(n540), .ZN(n521) );
  NAND2_X1 U623 ( .A1(n522), .A2(n521), .ZN(n637) );
  NAND2_X1 U624 ( .A1(n650), .A2(n637), .ZN(n536) );
  XOR2_X1 U625 ( .A(G122), .B(KEYINPUT7), .Z(n524) );
  XNOR2_X1 U626 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(n527), .ZN(n706) );
  NOR2_X1 U628 ( .A1(G902), .A2(n706), .ZN(n529) );
  XNOR2_X1 U629 ( .A(G478), .B(n529), .ZN(n548) );
  INV_X1 U630 ( .A(n548), .ZN(n534) );
  XOR2_X1 U631 ( .A(KEYINPUT13), .B(KEYINPUT104), .Z(n531) );
  XNOR2_X1 U632 ( .A(KEYINPUT103), .B(G475), .ZN(n530) );
  NOR2_X1 U633 ( .A1(G902), .A2(n532), .ZN(n533) );
  NAND2_X1 U634 ( .A1(n534), .A2(n549), .ZN(n651) );
  XNOR2_X1 U635 ( .A(KEYINPUT105), .B(n651), .ZN(n590) );
  NOR2_X1 U636 ( .A1(n611), .A2(n590), .ZN(n666) );
  INV_X1 U637 ( .A(n666), .ZN(n535) );
  NAND2_X1 U638 ( .A1(n536), .A2(n535), .ZN(n547) );
  XNOR2_X1 U639 ( .A(n537), .B(KEYINPUT107), .ZN(n538) );
  NAND2_X1 U640 ( .A1(n538), .A2(n347), .ZN(n539) );
  INV_X1 U641 ( .A(n540), .ZN(n541) );
  XNOR2_X1 U642 ( .A(KEYINPUT34), .B(KEYINPUT81), .ZN(n543) );
  NOR2_X1 U643 ( .A1(n549), .A2(n548), .ZN(n544) );
  XNOR2_X1 U644 ( .A(KEYINPUT108), .B(n544), .ZN(n599) );
  INV_X1 U645 ( .A(n664), .ZN(n552) );
  XNOR2_X1 U646 ( .A(KEYINPUT22), .B(KEYINPUT67), .ZN(n553) );
  XOR2_X1 U647 ( .A(n571), .B(KEYINPUT82), .Z(n555) );
  NOR2_X2 U648 ( .A1(n558), .A2(n409), .ZN(n563) );
  AND2_X1 U649 ( .A1(n559), .A2(n563), .ZN(n560) );
  NAND2_X1 U650 ( .A1(n560), .A2(n572), .ZN(n641) );
  NAND2_X1 U651 ( .A1(n565), .A2(KEYINPUT44), .ZN(n561) );
  NOR2_X1 U652 ( .A1(n572), .A2(n347), .ZN(n562) );
  NAND2_X1 U653 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U654 ( .A(KEYINPUT106), .B(n564), .ZN(n741) );
  NOR2_X1 U655 ( .A1(KEYINPUT44), .A2(n565), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n566), .A2(n407), .ZN(n567) );
  NAND2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U658 ( .A(n570), .ZN(n619) );
  INV_X1 U659 ( .A(n572), .ZN(n674) );
  NOR2_X1 U660 ( .A1(G900), .A2(n573), .ZN(n574) );
  NAND2_X1 U661 ( .A1(G953), .A2(n574), .ZN(n575) );
  XNOR2_X1 U662 ( .A(n575), .B(KEYINPUT110), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n673), .A2(n584), .ZN(n578) );
  XNOR2_X1 U665 ( .A(KEYINPUT72), .B(n579), .ZN(n592) );
  NOR2_X1 U666 ( .A1(n409), .A2(n605), .ZN(n580) );
  NAND2_X1 U667 ( .A1(n580), .A2(n661), .ZN(n581) );
  XNOR2_X1 U668 ( .A(n581), .B(KEYINPUT43), .ZN(n583) );
  BUF_X1 U669 ( .A(n582), .Z(n588) );
  INV_X1 U670 ( .A(n588), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n583), .A2(n602), .ZN(n657) );
  NAND2_X1 U672 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U673 ( .A(KEYINPUT38), .B(n588), .Z(n662) );
  NAND2_X1 U674 ( .A1(n600), .A2(n662), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n610), .A2(n590), .ZN(n656) );
  XOR2_X1 U676 ( .A(KEYINPUT111), .B(n591), .Z(n596) );
  XOR2_X1 U677 ( .A(KEYINPUT112), .B(KEYINPUT28), .Z(n594) );
  NAND2_X1 U678 ( .A1(n677), .A2(n592), .ZN(n593) );
  XNOR2_X1 U679 ( .A(n594), .B(n593), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n596), .A2(n595), .ZN(n613) );
  INV_X1 U681 ( .A(n613), .ZN(n598) );
  NAND2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n646) );
  NAND2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n645) );
  XOR2_X1 U685 ( .A(KEYINPUT83), .B(n645), .Z(n603) );
  NOR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT36), .B(KEYINPUT90), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n607), .B(n606), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n662), .A2(n661), .ZN(n665) );
  NOR2_X1 U690 ( .A1(n665), .A2(n664), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT41), .ZN(n691) );
  NOR2_X1 U692 ( .A1(n613), .A2(n691), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT42), .ZN(n738) );
  NOR2_X1 U694 ( .A1(n740), .A2(n738), .ZN(n616) );
  XNOR2_X1 U695 ( .A(KEYINPUT46), .B(KEYINPUT88), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n616), .B(n615), .ZN(n617) );
  XOR2_X1 U697 ( .A(n619), .B(KEYINPUT87), .Z(n620) );
  NAND2_X1 U698 ( .A1(n620), .A2(KEYINPUT2), .ZN(n621) );
  AND2_X1 U699 ( .A1(G472), .A2(n622), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n625), .B(KEYINPUT93), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n714), .A2(n630), .ZN(n633) );
  INV_X1 U703 ( .A(KEYINPUT63), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(G57) );
  NOR2_X1 U705 ( .A1(n648), .A2(n637), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n634), .B(KEYINPUT115), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(G6) );
  NOR2_X1 U708 ( .A1(n651), .A2(n637), .ZN(n639) );
  XNOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U711 ( .A(G107), .B(n640), .ZN(G9) );
  XNOR2_X1 U712 ( .A(n641), .B(G110), .ZN(G12) );
  NOR2_X1 U713 ( .A1(n651), .A2(n646), .ZN(n643) );
  XNOR2_X1 U714 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(G128), .B(n644), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n645), .Z(G45) );
  NOR2_X1 U718 ( .A1(n648), .A2(n646), .ZN(n647) );
  XOR2_X1 U719 ( .A(G146), .B(n647), .Z(G48) );
  NOR2_X1 U720 ( .A1(n648), .A2(n650), .ZN(n649) );
  XOR2_X1 U721 ( .A(G113), .B(n649), .Z(G15) );
  NOR2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U723 ( .A(G116), .B(n652), .Z(G18) );
  XOR2_X1 U724 ( .A(G125), .B(KEYINPUT37), .Z(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(G27) );
  XOR2_X1 U726 ( .A(G134), .B(KEYINPUT117), .Z(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(G36) );
  XNOR2_X1 U728 ( .A(G140), .B(n657), .ZN(G42) );
  XNOR2_X1 U729 ( .A(n658), .B(KEYINPUT2), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n659), .B(KEYINPUT86), .ZN(n695) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n660), .A2(n669), .ZN(n686) );
  NOR2_X1 U736 ( .A1(n671), .A2(n409), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT50), .B(n672), .Z(n680) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U740 ( .A1(n349), .A2(n676), .ZN(n678) );
  XNOR2_X1 U741 ( .A(KEYINPUT118), .B(n678), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(KEYINPUT51), .B(n683), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n684), .A2(n691), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U747 ( .A(n687), .B(KEYINPUT119), .Z(n688) );
  XNOR2_X1 U748 ( .A(KEYINPUT52), .B(n688), .ZN(n689) );
  NOR2_X1 U749 ( .A1(n690), .A2(n689), .ZN(n693) );
  NOR2_X1 U750 ( .A1(n660), .A2(n691), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n696), .A2(G953), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n697), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U755 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n699), .B(KEYINPUT57), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n708), .A2(G469), .ZN(n702) );
  XOR2_X1 U759 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U760 ( .A1(n714), .A2(n704), .ZN(G54) );
  NAND2_X1 U761 ( .A1(G478), .A2(n348), .ZN(n705) );
  XNOR2_X1 U762 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n714), .A2(n707), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n348), .A2(G217), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U766 ( .A(n380), .B(n715), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n718), .A2(n717), .ZN(n725) );
  NAND2_X1 U768 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n719), .B(KEYINPUT124), .ZN(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U771 ( .A1(G898), .A2(n721), .ZN(n723) );
  NAND2_X1 U772 ( .A1(n379), .A2(n731), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(G69) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(n729) );
  XOR2_X1 U776 ( .A(n728), .B(n729), .Z(n733) );
  XOR2_X1 U777 ( .A(n733), .B(n730), .Z(n732) );
  NAND2_X1 U778 ( .A1(n732), .A2(n731), .ZN(n737) );
  XNOR2_X1 U779 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n737), .A2(n736), .ZN(G72) );
  XNOR2_X1 U783 ( .A(G137), .B(KEYINPUT127), .ZN(n739) );
  XNOR2_X1 U784 ( .A(n739), .B(n738), .ZN(G39) );
  XOR2_X1 U785 ( .A(G131), .B(n740), .Z(G33) );
  XNOR2_X1 U786 ( .A(G101), .B(n741), .ZN(G3) );
  XNOR2_X1 U787 ( .A(G122), .B(KEYINPUT125), .ZN(n743) );
  XOR2_X1 U788 ( .A(n743), .B(n407), .Z(G24) );
  XNOR2_X1 U789 ( .A(G119), .B(KEYINPUT126), .ZN(n744) );
endmodule

