

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(KEYINPUT104), .ZN(n716) );
  NOR2_X1 U554 ( .A1(n975), .A2(n632), .ZN(n633) );
  XNOR2_X1 U555 ( .A(n695), .B(n694), .ZN(n718) );
  NAND2_X1 U556 ( .A1(n626), .A2(n625), .ZN(n687) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n626) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n521), .ZN(n882) );
  NOR2_X1 U559 ( .A1(G651), .A2(n579), .ZN(n787) );
  NOR2_X1 U560 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U561 ( .A1(n623), .A2(n622), .ZN(n975) );
  NOR2_X2 U562 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n519), .Z(n879) );
  AND2_X1 U565 ( .A1(n879), .A2(G138), .ZN(n527) );
  INV_X1 U566 ( .A(G2105), .ZN(n521) );
  AND2_X1 U567 ( .A1(n521), .A2(G2104), .ZN(n878) );
  NAND2_X1 U568 ( .A1(G102), .A2(n878), .ZN(n520) );
  XOR2_X1 U569 ( .A(KEYINPUT91), .B(n520), .Z(n525) );
  NAND2_X1 U570 ( .A1(G126), .A2(n882), .ZN(n523) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U572 ( .A1(G114), .A2(n884), .ZN(n522) );
  AND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U575 ( .A1(n527), .A2(n526), .ZN(G164) );
  NAND2_X1 U576 ( .A1(G101), .A2(n878), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(n528), .Z(n531) );
  NAND2_X1 U578 ( .A1(G125), .A2(n882), .ZN(n529) );
  XOR2_X1 U579 ( .A(n529), .B(KEYINPUT65), .Z(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U581 ( .A1(G137), .A2(n879), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G113), .A2(n884), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n579) );
  NAND2_X1 U585 ( .A1(n787), .A2(G52), .ZN(n538) );
  XOR2_X1 U586 ( .A(G651), .B(KEYINPUT66), .Z(n540) );
  NOR2_X1 U587 ( .A1(G543), .A2(n540), .ZN(n536) );
  XOR2_X2 U588 ( .A(KEYINPUT1), .B(n536), .Z(n788) );
  NAND2_X1 U589 ( .A1(G64), .A2(n788), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U591 ( .A(KEYINPUT68), .B(n539), .ZN(n546) );
  NOR2_X1 U592 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U593 ( .A1(n791), .A2(G90), .ZN(n542) );
  NOR2_X1 U594 ( .A1(n579), .A2(n540), .ZN(n792) );
  NAND2_X1 U595 ( .A1(G77), .A2(n792), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U597 ( .A(KEYINPUT9), .B(n543), .ZN(n544) );
  XNOR2_X1 U598 ( .A(KEYINPUT69), .B(n544), .ZN(n545) );
  NOR2_X1 U599 ( .A1(n546), .A2(n545), .ZN(G171) );
  NAND2_X1 U600 ( .A1(G89), .A2(n791), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT75), .B(n547), .Z(n548) );
  XNOR2_X1 U602 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G76), .A2(n792), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U605 ( .A(n551), .B(KEYINPUT5), .ZN(n556) );
  NAND2_X1 U606 ( .A1(n787), .A2(G51), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G63), .A2(n788), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n554), .Z(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U611 ( .A(n557), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(n787), .A2(G50), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G62), .A2(n788), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U616 ( .A1(n791), .A2(G88), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G75), .A2(n792), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U619 ( .A(KEYINPUT83), .B(n562), .Z(n563) );
  NOR2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U621 ( .A(KEYINPUT84), .B(n565), .Z(G303) );
  NAND2_X1 U622 ( .A1(n791), .A2(G86), .ZN(n566) );
  XOR2_X1 U623 ( .A(KEYINPUT81), .B(n566), .Z(n568) );
  NAND2_X1 U624 ( .A1(G61), .A2(n788), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U626 ( .A(KEYINPUT82), .B(n569), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G73), .A2(n792), .ZN(n570) );
  XOR2_X1 U628 ( .A(KEYINPUT2), .B(n570), .Z(n571) );
  NOR2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n787), .A2(G48), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(G305) );
  NAND2_X1 U632 ( .A1(G49), .A2(n787), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U635 ( .A1(n788), .A2(n577), .ZN(n578) );
  XNOR2_X1 U636 ( .A(n578), .B(KEYINPUT80), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G87), .A2(n579), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U639 ( .A1(n787), .A2(G47), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G60), .A2(n788), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U642 ( .A1(n791), .A2(G85), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G72), .A2(n792), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U645 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U646 ( .A(n588), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U647 ( .A1(G160), .A2(G40), .ZN(n624) );
  NOR2_X1 U648 ( .A1(n626), .A2(n624), .ZN(n747) );
  NAND2_X1 U649 ( .A1(G129), .A2(n882), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G117), .A2(n884), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U652 ( .A1(n878), .A2(G105), .ZN(n591) );
  XOR2_X1 U653 ( .A(KEYINPUT38), .B(n591), .Z(n592) );
  NOR2_X1 U654 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U655 ( .A1(n879), .A2(G141), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n595), .A2(n594), .ZN(n899) );
  AND2_X1 U657 ( .A1(n899), .A2(G1996), .ZN(n916) );
  NAND2_X1 U658 ( .A1(G119), .A2(n882), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G107), .A2(n884), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U661 ( .A1(G95), .A2(n878), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G131), .A2(n879), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U664 ( .A(KEYINPUT93), .B(n600), .Z(n601) );
  OR2_X1 U665 ( .A1(n602), .A2(n601), .ZN(n890) );
  AND2_X1 U666 ( .A1(n890), .A2(G1991), .ZN(n922) );
  OR2_X1 U667 ( .A1(n916), .A2(n922), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n747), .A2(n603), .ZN(n736) );
  XNOR2_X1 U669 ( .A(KEYINPUT92), .B(KEYINPUT34), .ZN(n607) );
  NAND2_X1 U670 ( .A1(G104), .A2(n878), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G140), .A2(n879), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n607), .B(n606), .ZN(n612) );
  NAND2_X1 U674 ( .A1(G128), .A2(n882), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G116), .A2(n884), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U677 ( .A(KEYINPUT35), .B(n610), .Z(n611) );
  NOR2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U679 ( .A(KEYINPUT36), .B(n613), .ZN(n891) );
  XNOR2_X1 U680 ( .A(G2067), .B(KEYINPUT37), .ZN(n745) );
  NOR2_X1 U681 ( .A1(n891), .A2(n745), .ZN(n913) );
  NAND2_X1 U682 ( .A1(n747), .A2(n913), .ZN(n743) );
  NAND2_X1 U683 ( .A1(n736), .A2(n743), .ZN(n733) );
  NAND2_X1 U684 ( .A1(n791), .A2(G81), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(KEYINPUT12), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G68), .A2(n792), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U688 ( .A(KEYINPUT13), .B(n617), .Z(n621) );
  NAND2_X1 U689 ( .A1(n788), .A2(G56), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(KEYINPUT14), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT71), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n787), .A2(G43), .ZN(n622) );
  INV_X1 U693 ( .A(n624), .ZN(n625) );
  INV_X1 U694 ( .A(G1996), .ZN(n627) );
  NOR2_X1 U695 ( .A1(n687), .A2(n627), .ZN(n629) );
  XNOR2_X1 U696 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(n631) );
  NAND2_X1 U698 ( .A1(n687), .A2(G1341), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U700 ( .A(KEYINPUT64), .B(n633), .Z(n648) );
  NAND2_X1 U701 ( .A1(n792), .A2(G79), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(KEYINPUT74), .ZN(n641) );
  NAND2_X1 U703 ( .A1(G92), .A2(n791), .ZN(n636) );
  NAND2_X1 U704 ( .A1(G54), .A2(n787), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U706 ( .A1(G66), .A2(n788), .ZN(n637) );
  XNOR2_X1 U707 ( .A(KEYINPUT73), .B(n637), .ZN(n638) );
  NOR2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U710 ( .A(KEYINPUT15), .B(n642), .Z(n985) );
  OR2_X1 U711 ( .A1(n648), .A2(n985), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(KEYINPUT98), .ZN(n647) );
  INV_X1 U713 ( .A(n687), .ZN(n670) );
  NOR2_X1 U714 ( .A1(n670), .A2(G1348), .ZN(n645) );
  NOR2_X1 U715 ( .A1(G2067), .A2(n687), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n648), .A2(n985), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n661) );
  NAND2_X1 U720 ( .A1(n670), .A2(G2072), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n651), .B(KEYINPUT27), .ZN(n653) );
  INV_X1 U722 ( .A(G1956), .ZN(n995) );
  NOR2_X1 U723 ( .A1(n995), .A2(n670), .ZN(n652) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n662) );
  NAND2_X1 U725 ( .A1(n787), .A2(G53), .ZN(n655) );
  NAND2_X1 U726 ( .A1(G65), .A2(n788), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n791), .A2(G91), .ZN(n657) );
  NAND2_X1 U729 ( .A1(G78), .A2(n792), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n972) );
  NAND2_X1 U732 ( .A1(n662), .A2(n972), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n662), .A2(n972), .ZN(n664) );
  XOR2_X1 U735 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n663) );
  XNOR2_X1 U736 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n668) );
  XNOR2_X1 U738 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n670), .A2(G1961), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n669), .B(KEYINPUT95), .ZN(n672) );
  XNOR2_X1 U742 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U743 ( .A1(n670), .A2(n944), .ZN(n671) );
  NAND2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n678), .A2(G171), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n685) );
  NAND2_X1 U747 ( .A1(G8), .A2(n687), .ZN(n729) );
  NOR2_X1 U748 ( .A1(G1966), .A2(n729), .ZN(n699) );
  NOR2_X1 U749 ( .A1(G2084), .A2(n687), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n699), .A2(n696), .ZN(n675) );
  NAND2_X1 U751 ( .A1(G8), .A2(n675), .ZN(n676) );
  XNOR2_X1 U752 ( .A(KEYINPUT30), .B(n676), .ZN(n677) );
  NOR2_X1 U753 ( .A1(G168), .A2(n677), .ZN(n681) );
  NOR2_X1 U754 ( .A1(G171), .A2(n678), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(KEYINPUT100), .ZN(n680) );
  NOR2_X1 U756 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U757 ( .A(n682), .B(KEYINPUT101), .ZN(n683) );
  XNOR2_X1 U758 ( .A(n683), .B(KEYINPUT31), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U760 ( .A(n686), .B(KEYINPUT102), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n697), .A2(G286), .ZN(n692) );
  NOR2_X1 U762 ( .A1(G1971), .A2(n729), .ZN(n689) );
  NOR2_X1 U763 ( .A1(G2090), .A2(n687), .ZN(n688) );
  NOR2_X1 U764 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U765 ( .A1(G303), .A2(n690), .ZN(n691) );
  NAND2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U767 ( .A1(n693), .A2(G8), .ZN(n695) );
  XOR2_X1 U768 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n694) );
  NAND2_X1 U769 ( .A1(G8), .A2(n696), .ZN(n701) );
  INV_X1 U770 ( .A(n697), .ZN(n698) );
  NOR2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n719) );
  XOR2_X1 U773 ( .A(G1981), .B(G305), .Z(n965) );
  INV_X1 U774 ( .A(n729), .ZN(n702) );
  NAND2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n978) );
  AND2_X1 U776 ( .A1(n702), .A2(n978), .ZN(n703) );
  NOR2_X1 U777 ( .A1(KEYINPUT33), .A2(n703), .ZN(n706) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NAND2_X1 U779 ( .A1(n969), .A2(KEYINPUT33), .ZN(n704) );
  NOR2_X1 U780 ( .A1(n704), .A2(n729), .ZN(n705) );
  NOR2_X1 U781 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U782 ( .A1(n965), .A2(n707), .ZN(n709) );
  AND2_X1 U783 ( .A1(n719), .A2(n709), .ZN(n708) );
  NAND2_X1 U784 ( .A1(n718), .A2(n708), .ZN(n715) );
  INV_X1 U785 ( .A(n709), .ZN(n713) );
  NOR2_X1 U786 ( .A1(G303), .A2(G1971), .ZN(n971) );
  NOR2_X1 U787 ( .A1(n969), .A2(n971), .ZN(n711) );
  INV_X1 U788 ( .A(KEYINPUT33), .ZN(n710) );
  AND2_X1 U789 ( .A1(n711), .A2(n710), .ZN(n712) );
  OR2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U792 ( .A(n717), .B(n716), .ZN(n725) );
  NAND2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n722) );
  NOR2_X1 U794 ( .A1(G2090), .A2(G303), .ZN(n720) );
  NAND2_X1 U795 ( .A1(G8), .A2(n720), .ZN(n721) );
  NAND2_X1 U796 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U797 ( .A1(n723), .A2(n729), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n731) );
  NOR2_X1 U799 ( .A1(G1981), .A2(G305), .ZN(n726) );
  XOR2_X1 U800 ( .A(n726), .B(KEYINPUT24), .Z(n727) );
  XNOR2_X1 U801 ( .A(KEYINPUT94), .B(n727), .ZN(n728) );
  NOR2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n735) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U806 ( .A1(n984), .A2(n747), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n750) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n899), .ZN(n932) );
  INV_X1 U809 ( .A(n736), .ZN(n739) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n890), .ZN(n918) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n918), .A2(n737), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n932), .A2(n740), .ZN(n741) );
  XOR2_X1 U815 ( .A(KEYINPUT39), .B(n741), .Z(n742) );
  XNOR2_X1 U816 ( .A(n742), .B(KEYINPUT105), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n891), .A2(n745), .ZN(n912) );
  NAND2_X1 U819 ( .A1(n746), .A2(n912), .ZN(n748) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U822 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U823 ( .A(G2443), .B(G2446), .Z(n753) );
  XNOR2_X1 U824 ( .A(G2427), .B(G2451), .ZN(n752) );
  XNOR2_X1 U825 ( .A(n753), .B(n752), .ZN(n759) );
  XOR2_X1 U826 ( .A(G2430), .B(G2454), .Z(n755) );
  XNOR2_X1 U827 ( .A(G1348), .B(G1341), .ZN(n754) );
  XNOR2_X1 U828 ( .A(n755), .B(n754), .ZN(n757) );
  XOR2_X1 U829 ( .A(G2435), .B(G2438), .Z(n756) );
  XNOR2_X1 U830 ( .A(n757), .B(n756), .ZN(n758) );
  XOR2_X1 U831 ( .A(n759), .B(n758), .Z(n760) );
  AND2_X1 U832 ( .A1(G14), .A2(n760), .ZN(G401) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G69), .ZN(G235) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U838 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U839 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n763) );
  INV_X1 U840 ( .A(G223), .ZN(n825) );
  NAND2_X1 U841 ( .A1(G567), .A2(n825), .ZN(n762) );
  XNOR2_X1 U842 ( .A(n763), .B(n762), .ZN(G234) );
  INV_X1 U843 ( .A(G860), .ZN(n833) );
  OR2_X1 U844 ( .A1(n975), .A2(n833), .ZN(G153) );
  INV_X1 U845 ( .A(G171), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G301), .A2(G868), .ZN(n764) );
  XNOR2_X1 U847 ( .A(n764), .B(KEYINPUT72), .ZN(n766) );
  INV_X1 U848 ( .A(G868), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n767), .A2(n985), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(G284) );
  INV_X1 U851 ( .A(n972), .ZN(G299) );
  NOR2_X1 U852 ( .A1(G286), .A2(n767), .ZN(n768) );
  XNOR2_X1 U853 ( .A(n768), .B(KEYINPUT76), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G299), .A2(G868), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n833), .A2(G559), .ZN(n771) );
  INV_X1 U857 ( .A(n985), .ZN(n859) );
  NAND2_X1 U858 ( .A1(n771), .A2(n859), .ZN(n772) );
  XNOR2_X1 U859 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n975), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n859), .A2(G868), .ZN(n773) );
  NOR2_X1 U862 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(G282) );
  NAND2_X1 U864 ( .A1(G99), .A2(n878), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G111), .A2(n884), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT78), .B(n778), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n882), .A2(G123), .ZN(n779) );
  XNOR2_X1 U869 ( .A(n779), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G135), .A2(n879), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U872 ( .A(KEYINPUT77), .B(n782), .Z(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n917) );
  XNOR2_X1 U874 ( .A(G2096), .B(n917), .ZN(n786) );
  INV_X1 U875 ( .A(G2100), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(G156) );
  NAND2_X1 U877 ( .A1(n787), .A2(G55), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G67), .A2(n788), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n791), .A2(G93), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U884 ( .A(n797), .B(KEYINPUT79), .Z(n834) );
  OR2_X1 U885 ( .A1(G868), .A2(n834), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT88), .ZN(n810) );
  XOR2_X1 U887 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n800) );
  XNOR2_X1 U888 ( .A(n972), .B(n834), .ZN(n799) );
  XNOR2_X1 U889 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U890 ( .A(KEYINPUT19), .B(n801), .ZN(n803) );
  XNOR2_X1 U891 ( .A(G305), .B(KEYINPUT85), .ZN(n802) );
  XNOR2_X1 U892 ( .A(n803), .B(n802), .ZN(n804) );
  XOR2_X1 U893 ( .A(n804), .B(G290), .Z(n805) );
  XNOR2_X1 U894 ( .A(G288), .B(n805), .ZN(n806) );
  XNOR2_X1 U895 ( .A(G303), .B(n806), .ZN(n855) );
  NAND2_X1 U896 ( .A1(G559), .A2(n859), .ZN(n807) );
  XOR2_X1 U897 ( .A(n975), .B(n807), .Z(n832) );
  XNOR2_X1 U898 ( .A(n855), .B(n832), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G868), .A2(n808), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n815), .Z(n816) );
  NOR2_X1 U909 ( .A1(G218), .A2(n816), .ZN(n817) );
  XOR2_X1 U910 ( .A(KEYINPUT89), .B(n817), .Z(n818) );
  NAND2_X1 U911 ( .A1(G96), .A2(n818), .ZN(n830) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n830), .ZN(n819) );
  XNOR2_X1 U913 ( .A(n819), .B(KEYINPUT90), .ZN(n823) );
  NAND2_X1 U914 ( .A1(G120), .A2(G108), .ZN(n820) );
  NOR2_X1 U915 ( .A1(G235), .A2(n820), .ZN(n821) );
  NAND2_X1 U916 ( .A1(G57), .A2(n821), .ZN(n831) );
  NAND2_X1 U917 ( .A1(G567), .A2(n831), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n906) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n906), .A2(n824), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U922 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U925 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U927 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XNOR2_X1 U929 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  NAND2_X1 U934 ( .A1(n833), .A2(n832), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(n834), .Z(G145) );
  XOR2_X1 U936 ( .A(KEYINPUT42), .B(G2090), .Z(n837) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n838), .B(G2096), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2678), .Z(n842) );
  XNOR2_X1 U943 ( .A(KEYINPUT109), .B(G2100), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(G227) );
  XNOR2_X1 U946 ( .A(G1981), .B(KEYINPUT41), .ZN(n854) );
  XOR2_X1 U947 ( .A(G1961), .B(G1956), .Z(n846) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1966), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U953 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U954 ( .A(G2474), .B(KEYINPUT110), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(G229) );
  XNOR2_X1 U957 ( .A(G286), .B(n855), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n975), .B(G171), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  NOR2_X1 U961 ( .A1(G37), .A2(n860), .ZN(G397) );
  NAND2_X1 U962 ( .A1(G124), .A2(n882), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G100), .A2(n878), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT111), .B(n862), .Z(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G136), .A2(n879), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G112), .A2(n884), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G130), .A2(n882), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G118), .A2(n884), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G106), .A2(n878), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G142), .A2(n879), .ZN(n871) );
  NAND2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U977 ( .A(KEYINPUT112), .B(n873), .Z(n874) );
  XNOR2_X1 U978 ( .A(KEYINPUT45), .B(n874), .ZN(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U980 ( .A(G160), .B(n877), .ZN(n895) );
  NAND2_X1 U981 ( .A1(G103), .A2(n878), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G139), .A2(n879), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n889) );
  NAND2_X1 U984 ( .A1(n882), .A2(G127), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n883), .B(KEYINPUT114), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G115), .A2(n884), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n925) );
  XNOR2_X1 U990 ( .A(n925), .B(n917), .ZN(n893) );
  XOR2_X1 U991 ( .A(n891), .B(n890), .Z(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n903) );
  XOR2_X1 U994 ( .A(KEYINPUT115), .B(KEYINPUT113), .Z(n897) );
  XNOR2_X1 U995 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n898), .B(G162), .Z(n901) );
  XOR2_X1 U998 ( .A(G164), .B(n899), .Z(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(n905), .ZN(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT108), .B(n906), .Z(G319) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n909) );
  AND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n911), .A2(G319), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G303), .ZN(G166) );
  INV_X1 U1012 ( .A(G57), .ZN(G237) );
  INV_X1 U1013 ( .A(n912), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n924) );
  XOR2_X1 U1015 ( .A(G160), .B(G2084), .Z(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n937) );
  XNOR2_X1 U1021 ( .A(G2072), .B(n925), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(G164), .B(G2078), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n926), .B(KEYINPUT118), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n929), .B(KEYINPUT119), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n930), .ZN(n935) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n961) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n961), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n956) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(G2072), .B(G33), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(KEYINPUT120), .B(n943), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(n944), .B(G27), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1043 ( .A(G32), .B(G1996), .Z(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT121), .B(n947), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(KEYINPUT122), .B(n950), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G25), .B(G1991), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n957), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n961), .B(n960), .ZN(n963) );
  INV_X1 U1056 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n964), .ZN(n1022) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT123), .ZN(n968) );
  XOR2_X1 U1063 ( .A(KEYINPUT57), .B(n968), .Z(n992) );
  XNOR2_X1 U1064 ( .A(KEYINPUT124), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n982) );
  XNOR2_X1 U1066 ( .A(n972), .B(G1956), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1341), .B(KEYINPUT125), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(G1961), .B(G301), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G1348), .B(n985), .Z(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT126), .B(n990), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n1020) );
  INV_X1 U1082 ( .A(G16), .ZN(n1018) );
  XNOR2_X1 U1083 ( .A(G20), .B(n995), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(G6), .B(G1981), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(KEYINPUT59), .B(G1348), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(G4), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n1003) );
  XNOR2_X1 U1092 ( .A(n1004), .B(n1003), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G5), .B(G1961), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(G1986), .B(G24), .Z(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

