//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G125), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT68), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(KEYINPUT3), .B2(new_n470), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n480));
  OAI211_X1 g055(.A(G137), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G101), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n466), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OAI21_X1  g061(.A(KEYINPUT69), .B1(new_n468), .B2(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(new_n469), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n488), .A2(new_n477), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n466), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT70), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  AND3_X1   g075(.A1(new_n466), .A2(G102), .A3(G2104), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n466), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT4), .A2(G138), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n488), .A2(new_n466), .A3(new_n477), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(G126), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n508));
  NAND2_X1  g083(.A1(G114), .A2(G2104), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n466), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(G164));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI211_X1 g088(.A(G50), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n516), .B(new_n518), .C1(new_n512), .C2(new_n513), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT71), .A2(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT71), .A2(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n514), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n516), .A2(new_n518), .A3(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT6), .B(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n516), .A2(new_n518), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n530), .B1(new_n532), .B2(new_n533), .C1(new_n534), .C2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  XNOR2_X1  g112(.A(KEYINPUT5), .B(G543), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n524), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n532), .A2(new_n541), .B1(new_n519), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n524), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT72), .B(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n532), .A2(new_n547), .B1(new_n519), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NOR2_X1   g131(.A1(new_n512), .A2(new_n513), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n515), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n558), .A2(KEYINPUT73), .A3(G53), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n532), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n562), .A3(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(new_n519), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n538), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n524), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n560), .B(new_n568), .C1(new_n532), .C2(new_n561), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n563), .A2(new_n565), .A3(new_n567), .A4(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  NAND4_X1  g146(.A1(new_n538), .A2(new_n531), .A3(new_n520), .A4(new_n521), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n538), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n514), .B(new_n572), .C1(new_n573), .C2(new_n524), .ZN(G303));
  NAND2_X1  g149(.A1(new_n564), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n558), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n538), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n524), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n535), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n584), .A2(KEYINPUT74), .A3(G651), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n581), .A2(new_n585), .B1(G48), .B2(new_n558), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n564), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n524), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n532), .A2(new_n591), .B1(new_n519), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n564), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n519), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n535), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n597), .A2(new_n600), .B1(G651), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n558), .A2(G54), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n596), .B1(new_n606), .B2(G868), .ZN(G321));
  XOR2_X1   g182(.A(G321), .B(KEYINPUT75), .Z(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND3_X1  g189(.A1(new_n606), .A2(KEYINPUT76), .A3(new_n613), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n604), .A2(new_n605), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G559), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n491), .A2(G123), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT77), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n494), .A2(G135), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NOR2_X1   g204(.A1(new_n470), .A2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n464), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2100), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n641), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT78), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT17), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n660), .C1(new_n658), .C2(new_n654), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT79), .ZN(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n665), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n671), .A3(new_n669), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(KEYINPUT20), .A3(new_n668), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n672), .B(new_n674), .C1(new_n676), .C2(new_n671), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT80), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(G19), .ZN(new_n685));
  OAI21_X1  g260(.A(KEYINPUT85), .B1(new_n685), .B2(G16), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n685), .A2(KEYINPUT85), .A3(G16), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n687), .C1(new_n550), .C2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G1341), .Z(new_n690));
  NAND4_X1  g265(.A1(new_n624), .A2(G29), .A3(new_n626), .A4(new_n627), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G11), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(G28), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n694), .B2(G28), .ZN(new_n696));
  NAND2_X1  g271(.A1(G171), .A2(G16), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G5), .B2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n690), .A2(new_n691), .A3(new_n692), .A4(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G34), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT24), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT24), .ZN(new_n704));
  AOI21_X1  g279(.A(G29), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n485), .B2(G29), .ZN(new_n706));
  INV_X1    g281(.A(G2084), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G168), .A2(new_n688), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n688), .B2(G21), .ZN(new_n710));
  INV_X1    g285(.A(G1966), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n708), .B1(new_n699), .B2(new_n698), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n693), .A2(G27), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G164), .B2(new_n693), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT93), .B(G2078), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR4_X1   g292(.A1(new_n701), .A2(new_n712), .A3(new_n713), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n693), .A2(G32), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n494), .A2(G141), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n491), .A2(G129), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n630), .A2(G105), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n720), .A2(new_n721), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n719), .B1(new_n726), .B2(new_n693), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n706), .A2(new_n707), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT91), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n688), .A2(G4), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n606), .B2(new_n688), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1348), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n688), .A2(G20), .ZN(new_n737));
  OAI211_X1 g312(.A(KEYINPUT23), .B(new_n737), .C1(new_n610), .C2(new_n688), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT23), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT95), .B(G1956), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n718), .A2(new_n730), .A3(new_n736), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n464), .A2(G127), .ZN(new_n743));
  INV_X1    g318(.A(G115), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n470), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G2105), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n489), .A2(G139), .A3(new_n466), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n630), .A2(G103), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n749), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n750), .B1(new_n749), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n693), .A2(G33), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT90), .ZN(new_n760));
  INV_X1    g335(.A(G2072), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n757), .A2(new_n762), .A3(new_n758), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n761), .B1(new_n760), .B2(new_n763), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n499), .A2(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n693), .A2(G35), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n767), .A3(new_n769), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(G2090), .ZN(new_n774));
  INV_X1    g349(.A(new_n772), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n766), .B(G2090), .C1(new_n775), .C2(new_n770), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n774), .A2(new_n777), .B1(G2090), .B2(new_n773), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n742), .A2(new_n764), .A3(new_n765), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n693), .A2(G26), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n494), .A2(G140), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT86), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT86), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n782), .A2(new_n783), .B1(G128), .B2(new_n491), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n780), .B1(new_n788), .B2(new_n693), .ZN(new_n789));
  MUX2_X1   g364(.A(new_n780), .B(new_n789), .S(KEYINPUT28), .Z(new_n790));
  INV_X1    g365(.A(G2067), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n688), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n688), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT83), .B(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n688), .B1(new_n586), .B2(new_n587), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT32), .B(G1981), .Z(new_n800));
  AND2_X1   g375(.A1(new_n688), .A2(G6), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT84), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n688), .A2(G23), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G288), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G1976), .ZN(new_n811));
  AOI211_X1 g386(.A(KEYINPUT33), .B(new_n806), .C1(G288), .C2(G16), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(G1976), .B1(new_n809), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n804), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n805), .B1(new_n804), .B2(new_n816), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n793), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n693), .A2(G25), .ZN(new_n821));
  INV_X1    g396(.A(G131), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n493), .A2(KEYINPUT81), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT81), .B1(new_n493), .B2(new_n822), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n823), .A2(new_n824), .B1(G119), .B2(new_n491), .ZN(new_n825));
  OR2_X1    g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT82), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n821), .B1(new_n830), .B2(new_n693), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n688), .A2(G24), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n594), .B2(new_n688), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(G1986), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n833), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n804), .A2(new_n816), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT84), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n840), .A2(KEYINPUT34), .A3(new_n817), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n836), .A2(G1986), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n820), .A2(new_n838), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n779), .B(new_n792), .C1(new_n844), .C2(new_n845), .ZN(G150));
  NAND2_X1  g421(.A1(G150), .A2(KEYINPUT96), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(KEYINPUT36), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n792), .A4(new_n779), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(G311));
  AOI22_X1  g426(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n524), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT97), .B(G55), .Z(new_n854));
  XOR2_X1   g429(.A(KEYINPUT98), .B(G93), .Z(new_n855));
  OAI22_X1  g430(.A1(new_n532), .A2(new_n854), .B1(new_n519), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n606), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  INV_X1    g436(.A(new_n550), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n853), .A2(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n550), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT39), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n861), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n859), .B1(new_n868), .B2(G860), .ZN(G145));
  XNOR2_X1  g444(.A(new_n628), .B(new_n829), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n485), .B(KEYINPUT99), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n499), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n870), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n756), .A2(G164), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n491), .A2(G130), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n494), .A2(G142), .ZN(new_n877));
  NOR2_X1   g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n725), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OAI221_X1 g457(.A(new_n746), .B1(new_n510), .B2(new_n507), .C1(new_n754), .C2(new_n755), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n875), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n875), .B2(new_n883), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n787), .B(new_n632), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n632), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n787), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n875), .A2(new_n883), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n881), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n892), .B2(new_n884), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n874), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n870), .B(new_n872), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n890), .A3(new_n884), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(new_n594), .B(KEYINPUT100), .ZN(new_n902));
  XNOR2_X1  g477(.A(G288), .B(G303), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G305), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n619), .B(new_n866), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n610), .A2(new_n606), .ZN(new_n912));
  NAND2_X1  g487(.A1(G299), .A2(new_n617), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(KEYINPUT41), .A3(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n864), .A2(new_n865), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n619), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n916), .B(new_n920), .C1(new_n908), .C2(new_n909), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT101), .A4(KEYINPUT42), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(G868), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n863), .A2(G868), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT102), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(G295));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n933), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n917), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n864), .B2(new_n865), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(G171), .B(G286), .Z(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n866), .A2(KEYINPUT103), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n915), .A2(new_n914), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n941), .A2(new_n944), .A3(new_n913), .A4(new_n912), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n908), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n947), .A2(new_n907), .A3(new_n906), .A4(new_n948), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n895), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n950), .A2(new_n951), .A3(new_n954), .A4(new_n895), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT44), .Z(G397));
  NAND2_X1  g532(.A1(G299), .A2(KEYINPUT114), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT57), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n507), .B2(new_n510), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT45), .B(new_n960), .C1(new_n507), .C2(new_n510), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n476), .A2(G40), .A3(new_n484), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT56), .B(G2072), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(new_n960), .C1(new_n507), .C2(new_n510), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1956), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n972), .A2(KEYINPUT113), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT113), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n959), .B(new_n968), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1348), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n979));
  INV_X1    g554(.A(new_n475), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n474), .B1(new_n473), .B2(G2105), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n484), .B(G40), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n961), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n979), .B1(new_n983), .B2(new_n791), .ZN(new_n984));
  NOR4_X1   g559(.A1(new_n982), .A2(new_n961), .A3(KEYINPUT115), .A4(G2067), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n978), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n976), .A2(new_n606), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n988));
  INV_X1    g563(.A(new_n959), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  INV_X1    g567(.A(new_n961), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n966), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT58), .B(G1341), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n966), .A2(new_n963), .A3(new_n997), .A4(new_n964), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n862), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n992), .B1(new_n1000), .B2(KEYINPUT59), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(KEYINPUT117), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n999), .B2(new_n1003), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT61), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n990), .A2(new_n1008), .A3(new_n976), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n990), .B2(new_n976), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n986), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n986), .A2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n606), .ZN(new_n1017));
  AOI211_X1 g592(.A(KEYINPUT118), .B(new_n617), .C1(new_n986), .C2(new_n1012), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n966), .A2(new_n993), .A3(new_n791), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT115), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n983), .A2(new_n979), .A3(new_n791), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT60), .B1(new_n1023), .B2(new_n978), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT118), .B1(new_n1024), .B2(new_n617), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1016), .A2(new_n1015), .A3(new_n606), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1013), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1019), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n991), .B1(new_n1011), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n966), .A2(new_n963), .A3(new_n964), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n711), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n966), .A2(new_n969), .A3(new_n707), .A4(new_n971), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(G168), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1034), .B2(G8), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT51), .B1(new_n1036), .B2(G168), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n972), .A2(new_n699), .ZN(new_n1042));
  INV_X1    g617(.A(G2078), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n966), .A2(new_n963), .A3(new_n1043), .A4(new_n964), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(KEYINPUT119), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT53), .B1(new_n1044), .B2(KEYINPUT119), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT120), .B(new_n1042), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(G171), .B(KEYINPUT54), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT55), .B(G8), .C1(new_n523), .C2(new_n527), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT105), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT105), .ZN(new_n1059));
  NAND4_X1  g634(.A1(G303), .A2(new_n1059), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT106), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(G166), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(new_n1060), .A3(KEYINPUT106), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT107), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT107), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1063), .A2(new_n1070), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1971), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1031), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2090), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n966), .A2(new_n969), .A3(new_n1075), .A4(new_n971), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1981), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n586), .A2(new_n1080), .A3(new_n587), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n531), .A2(G48), .A3(G543), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT108), .B(G86), .Z(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n519), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT109), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n584), .A2(G651), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1087), .C1(new_n519), .C2(new_n1083), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G1981), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n983), .A2(new_n1065), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1081), .A2(new_n1090), .A3(KEYINPUT49), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G288), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G1976), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n994), .A2(G8), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT52), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n811), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1096), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1069), .A2(new_n1077), .A3(G8), .A4(new_n1071), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1079), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1050), .B1(new_n473), .B2(G2105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n484), .A2(G40), .A3(new_n1043), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n965), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(new_n1051), .A3(new_n1042), .A4(new_n1054), .ZN(new_n1109));
  AND4_X1   g684(.A1(new_n1041), .A2(new_n1056), .A3(new_n1105), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1029), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1079), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1040), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(KEYINPUT121), .A3(G171), .A4(new_n1053), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1035), .ZN(new_n1116));
  AOI21_X1  g691(.A(G168), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1117));
  OAI211_X1 g692(.A(G8), .B(new_n1034), .C1(new_n1117), .C2(new_n1030), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1118), .A3(new_n1113), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1105), .A2(new_n1119), .A3(new_n1053), .A4(G171), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1041), .A2(KEYINPUT62), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1096), .A2(new_n811), .A3(new_n1097), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1081), .B(KEYINPUT110), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT111), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT111), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1129), .A3(new_n1126), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1094), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1103), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1104), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT63), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1105), .A2(G168), .A3(new_n1039), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1112), .A2(new_n1038), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(new_n1134), .A3(KEYINPUT63), .A4(G168), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1111), .A2(new_n1124), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n963), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n966), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n784), .A2(new_n791), .A3(new_n786), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n791), .B1(new_n784), .B2(new_n786), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n725), .A2(G1996), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1145), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1144), .A2(G1996), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT104), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n726), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n829), .A2(new_n832), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n829), .A2(new_n832), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1145), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1151), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1144), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1142), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1154), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1144), .B1(new_n1166), .B2(new_n1149), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1156), .B(KEYINPUT122), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1164), .B1(new_n1169), .B2(new_n1146), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1146), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT123), .B(new_n1171), .C1(new_n1172), .C2(new_n1168), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1173), .A3(new_n1145), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1158), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1151), .A2(KEYINPUT125), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1144), .A2(new_n1159), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1145), .B1(new_n1148), .B2(new_n725), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT124), .B(KEYINPUT46), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1153), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1153), .B1(new_n1185), .B2(KEYINPUT46), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1182), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT47), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1174), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1163), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g765(.A1(new_n956), .A2(new_n649), .ZN(new_n1192));
  OR3_X1    g766(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1193));
  INV_X1    g767(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n900), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g769(.A(KEYINPUT127), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g770(.A(new_n649), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n953), .B2(new_n955), .ZN(new_n1198));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n1199));
  NAND4_X1  g773(.A1(new_n1198), .A2(new_n1199), .A3(new_n900), .A4(new_n1194), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1196), .A2(new_n1200), .ZN(G308));
  NAND3_X1  g775(.A1(new_n1198), .A2(new_n900), .A3(new_n1194), .ZN(G225));
endmodule


