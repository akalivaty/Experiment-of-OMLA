//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT18), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT89), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n210), .B1(new_n213), .B2(KEYINPUT88), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(G1gat), .B2(new_n211), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n214), .B(new_n215), .Z(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G43gat), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  INV_X1    g023(.A(G29gat), .ZN(new_n225));
  INV_X1    g024(.A(G36gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT84), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n225), .A2(new_n226), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT84), .B1(new_n227), .B2(new_n228), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n235));
  NOR3_X1   g034(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n221), .A2(new_n222), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n227), .A2(KEYINPUT85), .A3(new_n228), .ZN(new_n238));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n230), .B1(new_n239), .B2(KEYINPUT15), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(KEYINPUT17), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n216), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n234), .A2(new_n245), .A3(new_n241), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n234), .B2(new_n241), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT87), .B(new_n244), .C1(new_n246), .C2(new_n247), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G229gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n241), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT86), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n245), .A3(new_n241), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(new_n216), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n252), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n208), .A2(KEYINPUT89), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n209), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n243), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT87), .B1(new_n258), .B2(new_n244), .ZN(new_n265));
  INV_X1    g064(.A(new_n251), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n259), .A2(new_n216), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n209), .A3(new_n253), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(new_n216), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n253), .B(KEYINPUT13), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n207), .B1(new_n263), .B2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n267), .A2(new_n262), .A3(new_n253), .A4(new_n268), .ZN(new_n277));
  INV_X1    g076(.A(new_n209), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n279), .A2(new_n274), .A3(new_n269), .A4(new_n206), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT35), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n284));
  XNOR2_X1  g083(.A(G155gat), .B(G162gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n287));
  XNOR2_X1  g086(.A(G141gat), .B(G148gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(KEYINPUT72), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(KEYINPUT72), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(KEYINPUT74), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G141gat), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n285), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT75), .B(G162gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G162gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n309), .A3(G155gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT2), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT76), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  AND4_X1   g112(.A1(new_n284), .A2(new_n293), .A3(new_n294), .A4(new_n313), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n291), .A2(new_n292), .B1(new_n305), .B2(new_n312), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n284), .B1(new_n315), .B2(new_n294), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n293), .A2(new_n294), .A3(new_n313), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT79), .B1(new_n318), .B2(KEYINPUT3), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n315), .A2(new_n320), .A3(new_n321), .A4(new_n294), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G134gat), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n327));
  INV_X1    g126(.A(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G127gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT1), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT67), .B(G113gat), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n333), .A2(new_n325), .A3(new_n329), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n330), .A2(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT78), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n323), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n338), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n318), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n315), .A2(new_n294), .A3(new_n338), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n353), .A3(new_n344), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT80), .B1(new_n346), .B2(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n347), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n341), .A2(new_n356), .A3(new_n349), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n318), .A2(KEYINPUT77), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n315), .A2(new_n284), .A3(new_n294), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n343), .B1(new_n360), .B2(new_n340), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT5), .B1(new_n361), .B2(new_n349), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364));
  INV_X1    g163(.A(G85gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n370), .B(new_n352), .C1(new_n357), .C2(new_n362), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n314), .A2(new_n316), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n346), .B1(new_n375), .B2(new_n339), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(new_n350), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n341), .A2(new_n356), .A3(new_n349), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n346), .B(new_n344), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n339), .B1(new_n360), .B2(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n323), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n377), .A2(new_n378), .B1(new_n381), .B2(new_n351), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n368), .B(KEYINPUT82), .Z(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n369), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT65), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  AND2_X1   g195(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT28), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n399), .A2(KEYINPUT28), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n393), .A2(new_n395), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT64), .B1(new_n406), .B2(KEYINPUT24), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT64), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n388), .A2(KEYINPUT23), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(G169gat), .B2(G176gat), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n412), .A2(new_n414), .A3(new_n387), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(KEYINPUT25), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n403), .A2(new_n408), .A3(new_n404), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(new_n414), .A3(new_n387), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n402), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G197gat), .B(G204gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n428));
  AND2_X1   g227(.A1(G211gat), .A2(G218gat), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(G211gat), .A2(G218gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n430), .B(new_n432), .Z(new_n433));
  NAND2_X1  g232(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n433), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n424), .B(new_n435), .C1(new_n423), .C2(new_n425), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n434), .A2(KEYINPUT30), .A3(new_n442), .A4(new_n436), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n434), .A2(new_n442), .A3(new_n436), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT71), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n441), .B(new_n443), .C1(new_n445), .C2(KEYINPUT30), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n385), .A2(KEYINPUT83), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT29), .B1(new_n319), .B2(new_n322), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(new_n435), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT29), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT3), .B1(new_n435), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n294), .B2(new_n315), .ZN(new_n453));
  INV_X1    g252(.A(G228gat), .ZN(new_n454));
  INV_X1    g253(.A(G233gat), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n450), .A2(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  OAI221_X1 g256(.A(new_n457), .B1(new_n375), .B2(new_n452), .C1(new_n449), .C2(new_n435), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G50gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n458), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n422), .A2(new_n342), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n402), .A2(new_n421), .A3(new_n338), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(G227gat), .A2(G233gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n402), .A2(new_n421), .A3(new_n338), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n338), .B1(new_n402), .B2(new_n421), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n471), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT32), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT34), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n476), .B2(new_n480), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n474), .A2(new_n475), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G43gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G71gat), .B(G99gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n488), .A2(new_n489), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT68), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT33), .B1(new_n497), .B2(new_n479), .ZN(new_n498));
  INV_X1    g297(.A(new_n493), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n479), .ZN(new_n501));
  INV_X1    g300(.A(new_n484), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n502), .ZN(new_n503));
  AND4_X1   g302(.A1(new_n485), .A2(new_n494), .A3(new_n500), .A4(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n494), .A2(new_n500), .B1(new_n485), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n470), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n448), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n371), .B(new_n372), .C1(new_n382), .C2(new_n383), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n446), .B1(new_n509), .B2(new_n369), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(KEYINPUT83), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n283), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n504), .B2(new_n505), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n467), .A2(new_n469), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n490), .B1(new_n487), .B2(new_n493), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n498), .A2(new_n495), .A3(new_n499), .ZN(new_n517));
  INV_X1    g316(.A(new_n503), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n502), .B1(new_n501), .B2(KEYINPUT32), .ZN(new_n519));
  OAI22_X1  g318(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n494), .A2(new_n500), .A3(new_n485), .A4(new_n503), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT36), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n470), .B(KEYINPUT35), .C1(new_n504), .C2(new_n505), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n363), .A2(new_n368), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n372), .A3(new_n371), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n446), .B1(new_n527), .B2(new_n369), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT36), .B1(new_n520), .B2(new_n521), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n515), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n437), .A2(KEYINPUT37), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n434), .A2(new_n533), .A3(new_n436), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n440), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n532), .A2(KEYINPUT38), .A3(new_n440), .A4(new_n534), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n445), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n509), .A2(new_n369), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT39), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n361), .B2(new_n349), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n381), .B2(new_n349), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n341), .A2(new_n348), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n541), .A3(new_n350), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n383), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT40), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n383), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n363), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT40), .A4(new_n383), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n446), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n540), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n525), .A2(new_n528), .B1(new_n531), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n282), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(G71gat), .ZN(new_n558));
  INV_X1    g357(.A(G78gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n557), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  INV_X1    g364(.A(G64gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G57gat), .ZN(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G64gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT90), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n563), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n216), .B1(new_n556), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT20), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n556), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(G183gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G211gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n579), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G190gat), .B(G218gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n588));
  NOR2_X1   g387(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n588), .A2(new_n589), .B1(new_n365), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT7), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n365), .B2(new_n590), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n591), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n591), .A2(new_n597), .A3(new_n601), .A4(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n242), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n250), .B2(new_n251), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT41), .ZN(new_n608));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT92), .ZN(new_n610));
  OAI22_X1  g409(.A1(new_n259), .A2(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n587), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(KEYINPUT95), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n608), .ZN(new_n614));
  XOR2_X1   g413(.A(G134gat), .B(G162gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(KEYINPUT95), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n607), .A2(new_n611), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n586), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n623), .B2(new_n612), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n621), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n618), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n585), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT97), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n572), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n561), .A2(KEYINPUT90), .B1(new_n557), .B2(new_n564), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n567), .A2(new_n569), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT9), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n560), .A2(new_n557), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n632), .A2(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n604), .A2(KEYINPUT96), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n605), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n604), .B(new_n603), .C1(new_n573), .C2(KEYINPUT96), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n605), .A2(new_n642), .A3(new_n573), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n631), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n640), .A3(new_n630), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n628), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n555), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n527), .A2(new_n369), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n654), .A2(new_n447), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n660), .B2(new_n210), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT98), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G8gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  MUX2_X1   g463(.A(KEYINPUT42), .B(new_n661), .S(new_n664), .Z(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n514), .A2(new_n522), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n654), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n504), .A2(new_n505), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n669), .B1(new_n666), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n470), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n585), .ZN(new_n677));
  INV_X1    g476(.A(new_n624), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n617), .A2(new_n616), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n678), .A2(new_n625), .B1(new_n679), .B2(new_n613), .ZN(new_n680));
  INV_X1    g479(.A(new_n652), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT99), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n555), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n657), .A2(new_n225), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT100), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n686), .A2(KEYINPUT45), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n681), .A2(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n681), .A2(KEYINPUT101), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n282), .A3(new_n585), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n512), .A2(new_n554), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n680), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI211_X1 g497(.A(KEYINPUT44), .B(new_n627), .C1(new_n512), .C2(new_n554), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n694), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n225), .B1(new_n701), .B2(new_n657), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT45), .B1(new_n686), .B2(new_n687), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n688), .A2(new_n702), .A3(new_n703), .ZN(G1328gat));
  NOR3_X1   g503(.A1(new_n684), .A2(G36gat), .A3(new_n447), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  AOI21_X1  g505(.A(new_n226), .B1(new_n701), .B2(new_n446), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  OAI211_X1 g507(.A(new_n667), .B(new_n693), .C1(new_n697), .C2(new_n699), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT47), .B1(new_n710), .B2(KEYINPUT102), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n671), .A2(new_n219), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n684), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(new_n713), .ZN(G1330gat));
  AOI21_X1  g513(.A(new_n217), .B1(new_n701), .B2(new_n515), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n515), .A2(new_n217), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n684), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT48), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OR3_X1    g519(.A1(new_n715), .A2(new_n720), .A3(new_n717), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n715), .B2(new_n717), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n628), .A2(new_n281), .A3(new_n691), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n696), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  AOI211_X1 g526(.A(KEYINPUT104), .B(new_n727), .C1(new_n512), .C2(new_n554), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n656), .B(KEYINPUT105), .Z(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g531(.A(new_n447), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n735), .B(new_n736), .Z(G1333gat));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n729), .B2(new_n671), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n525), .A2(new_n528), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n531), .A2(new_n553), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n506), .B1(new_n510), .B2(KEYINPUT83), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n385), .A2(new_n447), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT83), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT35), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n725), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n696), .A2(new_n724), .A3(new_n725), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n750), .A2(new_n751), .A3(new_n739), .A4(new_n671), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n558), .B1(new_n740), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n558), .B1(new_n729), .B2(new_n667), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n738), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n750), .A2(new_n751), .A3(new_n671), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT107), .ZN(new_n759));
  AOI21_X1  g558(.A(G71gat), .B1(new_n759), .B2(new_n752), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(KEYINPUT50), .A3(new_n755), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n757), .A2(new_n761), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n729), .A2(new_n515), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g563(.A1(new_n677), .A2(new_n282), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n652), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n697), .B2(new_n699), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n656), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n696), .A2(new_n680), .A3(new_n766), .ZN(new_n771));
  NAND2_X1  g570(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n696), .A2(new_n680), .A3(new_n766), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n657), .A2(new_n365), .A3(new_n652), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n770), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n769), .B2(new_n447), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n771), .A2(new_n785), .A3(KEYINPUT51), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n771), .B2(new_n785), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n691), .A2(new_n447), .A3(G92gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(new_n777), .B2(new_n788), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(new_n783), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n792), .B2(new_n783), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n769), .B2(new_n668), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n670), .A2(G99gat), .A3(new_n681), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n778), .B2(new_n798), .ZN(G1338gat));
  OAI211_X1 g598(.A(new_n515), .B(new_n768), .C1(new_n697), .C2(new_n699), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n800), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n800), .B2(G106gat), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n691), .A2(G106gat), .A3(new_n470), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n786), .A2(new_n787), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n800), .A2(G106gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n778), .B2(new_n803), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n639), .A2(new_n640), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n642), .ZN(new_n811));
  INV_X1    g610(.A(new_n643), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n630), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n644), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n815), .B(new_n631), .C1(new_n641), .C2(new_n643), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n649), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n650), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n816), .A2(new_n649), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n819), .B2(new_n814), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n818), .B2(new_n820), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n822), .A2(new_n824), .B1(new_n276), .B2(new_n280), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n271), .A2(new_n273), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n253), .B1(new_n267), .B2(new_n268), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n205), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n280), .A2(new_n652), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n627), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n822), .A2(new_n824), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n280), .A2(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n680), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n677), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n628), .A2(new_n281), .A3(new_n652), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n506), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n657), .A2(new_n447), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n282), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n730), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n447), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n282), .A2(new_n335), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n841), .B2(new_n691), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n652), .A2(new_n332), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT116), .Z(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n846), .B2(new_n851), .ZN(G1341gat));
  OAI21_X1  g651(.A(G127gat), .B1(new_n841), .B2(new_n677), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n677), .A2(G127gat), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n853), .C1(new_n846), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1342gat));
  NAND2_X1  g659(.A1(new_n680), .A2(new_n328), .ZN(new_n861));
  OR3_X1    g660(.A1(new_n846), .A2(KEYINPUT56), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n841), .B2(new_n627), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT56), .B1(new_n846), .B2(new_n861), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n835), .A2(new_n837), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n515), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n667), .A2(new_n656), .A3(new_n446), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT118), .B1(new_n818), .B2(new_n820), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n819), .A2(new_n814), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n873), .A2(new_n874), .A3(new_n650), .A4(new_n817), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n829), .B1(new_n281), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n833), .B1(new_n877), .B2(new_n680), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n677), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n470), .B1(new_n879), .B2(new_n837), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n868), .B(new_n869), .C1(new_n867), .C2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G141gat), .B1(new_n881), .B2(new_n282), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT58), .B1(new_n882), .B2(KEYINPUT119), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n730), .A2(new_n447), .A3(new_n668), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n515), .A3(new_n866), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n282), .A2(G141gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n882), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  OAI221_X1 g689(.A(new_n882), .B1(KEYINPUT119), .B2(KEYINPUT58), .C1(new_n886), .C2(new_n888), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n881), .A2(new_n681), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .A3(new_n295), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n263), .A2(new_n275), .A3(new_n207), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n272), .B1(new_n268), .B2(new_n270), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n261), .B2(new_n209), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n206), .B1(new_n899), .B2(new_n279), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n870), .B(new_n875), .C1(new_n897), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n280), .A2(new_n652), .A3(new_n828), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n680), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n680), .A2(new_n821), .A3(new_n832), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n677), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n470), .B1(new_n905), .B2(new_n837), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n896), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n680), .A2(new_n821), .A3(new_n832), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n877), .B2(new_n680), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n836), .B1(new_n909), .B2(new_n677), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT120), .B(new_n867), .C1(new_n910), .C2(new_n470), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n585), .B1(new_n830), .B2(new_n833), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT57), .B(new_n515), .C1(new_n912), .C2(new_n836), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n907), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n652), .A3(new_n869), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n895), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n652), .A2(new_n295), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n894), .A2(new_n916), .B1(new_n886), .B2(new_n917), .ZN(G1345gat));
  NOR2_X1   g717(.A1(new_n886), .A2(new_n677), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n585), .A2(G155gat), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n919), .A2(G155gat), .B1(new_n881), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(new_n302), .B1(new_n881), .B2(new_n627), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n627), .A2(new_n302), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n886), .B2(new_n924), .ZN(G1347gat));
  INV_X1    g724(.A(new_n730), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n838), .A2(new_n446), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n282), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n657), .A2(new_n447), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n866), .A2(new_n507), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n282), .A2(G169gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT121), .Z(G1348gat));
  NAND2_X1  g732(.A1(new_n692), .A2(G176gat), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  INV_X1    g737(.A(G176gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n930), .B2(new_n681), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n936), .B(new_n937), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(new_n938), .B2(new_n940), .ZN(G1349gat));
  OAI21_X1  g741(.A(G183gat), .B1(new_n927), .B2(new_n677), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n585), .B1(new_n398), .B2(new_n397), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n930), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n927), .B2(new_n627), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n680), .A2(new_n396), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n930), .B2(new_n949), .ZN(G1351gat));
  XNOR2_X1  g749(.A(KEYINPUT124), .B(G197gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n730), .A2(new_n447), .A3(new_n667), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n914), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n282), .ZN(new_n954));
  INV_X1    g753(.A(new_n523), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n866), .A2(new_n955), .A3(new_n929), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n282), .A2(new_n951), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n953), .B2(new_n691), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n681), .A2(G204gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OR4_X1    g762(.A1(KEYINPUT125), .A2(new_n956), .A3(KEYINPUT62), .A4(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n956), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n966), .A3(new_n962), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT62), .B1(new_n956), .B2(new_n963), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n959), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n972), .A2(KEYINPUT126), .A3(new_n960), .A4(new_n964), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1353gat));
  OR3_X1    g773(.A1(new_n956), .A2(G211gat), .A3(new_n677), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n914), .A2(new_n585), .A3(new_n952), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(G211gat), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT63), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(KEYINPUT127), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT127), .B1(new_n977), .B2(new_n978), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  NAND2_X1  g782(.A1(new_n680), .A2(G218gat), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n953), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(G218gat), .B1(new_n965), .B2(new_n680), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


