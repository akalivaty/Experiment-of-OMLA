//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n192), .A2(KEYINPUT78), .A3(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT78), .B1(new_n192), .B2(new_n193), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n187), .A2(KEYINPUT79), .A3(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n187), .A2(G119), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(new_n199), .C1(new_n200), .C2(new_n193), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n195), .A3(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT68), .B(G128), .ZN(new_n203));
  OR3_X1    g017(.A1(new_n203), .A2(KEYINPUT76), .A3(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n192), .A2(KEYINPUT76), .ZN(new_n205));
  INV_X1    g019(.A(new_n200), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT24), .B(G110), .Z(new_n208));
  OAI22_X1  g022(.A1(new_n202), .A2(G110), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(G146), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(G110), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n207), .A2(KEYINPUT77), .A3(new_n208), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n215), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n214), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n208), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT77), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n219), .A2(new_n220), .A3(new_n223), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  INV_X1    g043(.A(G221), .ZN(new_n230));
  INV_X1    g044(.A(G234), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n230), .A2(new_n231), .A3(G953), .ZN(new_n232));
  XOR2_X1   g046(.A(new_n229), .B(new_n232), .Z(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT74), .B(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(new_n227), .A3(new_n233), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT25), .ZN(new_n240));
  OAI21_X1  g054(.A(G217), .B1(new_n236), .B2(new_n231), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n241), .B(KEYINPUT75), .Z(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n235), .A2(new_n243), .A3(new_n237), .A4(new_n238), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT80), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n240), .A2(new_n247), .A3(new_n242), .A4(new_n244), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n235), .A2(new_n238), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n242), .A2(G902), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G472), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  XNOR2_X1  g070(.A(G116), .B(G119), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT65), .A2(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT65), .A2(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(G146), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n261), .A2(KEYINPUT0), .A3(G128), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT0), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n187), .A3(KEYINPUT64), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(KEYINPUT0), .B2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n259), .A2(new_n260), .A3(G146), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n215), .A2(G143), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n266), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G137), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT11), .A2(G134), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT11), .A2(G134), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(G137), .B2(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n275), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n277), .B2(new_n279), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(G137), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT11), .A2(G134), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n287), .A2(new_n290), .A3(G131), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n265), .B(new_n274), .C1(new_n286), .C2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT66), .B(G137), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n285), .B(new_n275), .C1(new_n281), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g109(.A1(G134), .A2(G137), .ZN(new_n296));
  OAI211_X1 g110(.A(G131), .B(new_n296), .C1(new_n293), .C2(G134), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT1), .B1(new_n262), .B2(G146), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n188), .A3(new_n190), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n272), .B2(new_n273), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n261), .A2(new_n302), .A3(G128), .A4(new_n264), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n295), .B1(new_n294), .B2(new_n297), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n258), .B(new_n292), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n294), .A2(new_n297), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT69), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n304), .A3(new_n298), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n258), .A4(new_n292), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n304), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT67), .B1(new_n294), .B2(new_n297), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n292), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n258), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT26), .B(G101), .Z(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G210), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n322), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n331), .B(new_n292), .C1(new_n316), .C2(new_n317), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n311), .B2(new_n292), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n319), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n307), .A2(new_n328), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n292), .B1(new_n305), .B2(new_n306), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT30), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n258), .B1(new_n341), .B2(new_n332), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT31), .B1(new_n342), .B2(new_n337), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n330), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n330), .A2(new_n339), .A3(new_n343), .A4(KEYINPUT71), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n255), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT72), .B1(new_n348), .B2(KEYINPUT32), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n258), .B1(new_n311), .B2(new_n292), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n308), .B2(new_n313), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT29), .A3(new_n328), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n358), .B(KEYINPUT73), .Z(new_n359));
  INV_X1    g173(.A(new_n307), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n342), .A2(new_n360), .A3(new_n328), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n328), .B2(new_n321), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n359), .B(new_n237), .C1(KEYINPUT29), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G472), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n252), .B1(new_n355), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(G104), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT83), .B(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G104), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n368), .A2(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n369), .B2(new_n368), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT82), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G104), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n379), .A3(new_n368), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n378), .A2(G104), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n376), .A2(KEYINPUT82), .ZN(new_n384));
  OAI21_X1  g198(.A(G107), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G107), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n368), .A2(KEYINPUT83), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n381), .A2(new_n382), .A3(new_n385), .A4(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n375), .A2(KEYINPUT84), .A3(KEYINPUT4), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(G101), .C1(new_n373), .C2(new_n374), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n319), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n368), .A2(KEYINPUT83), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n387), .A2(G107), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n376), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n380), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G101), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n391), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n257), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n256), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G113), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n197), .A2(G116), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n409), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n401), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(G110), .B(G122), .Z(new_n418));
  OAI21_X1  g232(.A(new_n367), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n399), .B1(new_n394), .B2(new_n395), .ZN(new_n420));
  INV_X1    g234(.A(new_n416), .ZN(new_n421));
  NOR4_X1   g235(.A1(new_n420), .A2(new_n367), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n274), .A2(G125), .A3(new_n265), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(new_n212), .B2(new_n304), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(KEYINPUT90), .B2(KEYINPUT7), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n324), .A2(G224), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT89), .Z(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT7), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n427), .A2(new_n431), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n414), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n407), .B1(new_n409), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n418), .B(KEYINPUT8), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n391), .A2(new_n406), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n415), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n432), .A2(new_n433), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(G902), .B1(new_n424), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n421), .B1(new_n396), .B2(new_n400), .ZN(new_n445));
  INV_X1    g259(.A(new_n418), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT88), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT6), .B1(new_n447), .B2(new_n422), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n417), .A2(new_n418), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n426), .B(new_n429), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n442), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT91), .Z(new_n454));
  AOI21_X1  g268(.A(new_n366), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n454), .ZN(new_n456));
  INV_X1    g270(.A(new_n454), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n442), .B(new_n457), .C1(new_n450), .C2(new_n451), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n455), .B1(new_n459), .B2(new_n366), .ZN(new_n460));
  OAI21_X1  g274(.A(G214), .B1(G237), .B2(G902), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT86), .Z(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT9), .B(G234), .Z(new_n464));
  AOI21_X1  g278(.A(new_n230), .B1(new_n464), .B2(new_n254), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n286), .A2(new_n291), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n398), .A2(new_n265), .A3(new_n274), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n394), .B2(new_n395), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT10), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n262), .ZN(new_n472));
  NAND2_X1  g286(.A1(KEYINPUT65), .A2(G143), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n215), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n187), .B1(new_n474), .B2(KEYINPUT1), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n263), .B1(new_n476), .B2(G146), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n303), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n470), .B1(new_n479), .B2(new_n439), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n391), .A4(new_n406), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n467), .B1(new_n469), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n324), .A2(G227), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT81), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G140), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n488));
  INV_X1    g302(.A(new_n468), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n482), .B1(new_n396), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n490), .B2(new_n466), .ZN(new_n491));
  NOR4_X1   g305(.A1(new_n469), .A2(new_n482), .A3(KEYINPUT85), .A4(new_n467), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n483), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n407), .A2(new_n304), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n479), .A2(new_n439), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n467), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT12), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n396), .A2(new_n489), .ZN(new_n498));
  INV_X1    g312(.A(new_n482), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n466), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n488), .A3(new_n466), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n493), .B(G469), .C1(new_n503), .C2(new_n487), .ZN(new_n504));
  NAND2_X1  g318(.A1(G469), .A2(G902), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n483), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n508), .A2(new_n487), .B1(new_n509), .B2(new_n497), .ZN(new_n510));
  INV_X1    g324(.A(G469), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n237), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n465), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n259), .A2(new_n260), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n187), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n203), .A2(new_n262), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT96), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n191), .A2(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n476), .A2(G128), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(G134), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT97), .ZN(new_n524));
  XNOR2_X1  g338(.A(G116), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n370), .B(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  OR3_X1    g341(.A1(new_n515), .A2(new_n527), .A3(KEYINPUT13), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n515), .B2(KEYINPUT13), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n516), .B1(new_n515), .B2(KEYINPUT13), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n531), .B2(G134), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n522), .B2(G134), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n525), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n370), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n538));
  INV_X1    g352(.A(G122), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G116), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n368), .B1(new_n540), .B2(KEYINPUT14), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n522), .A2(G134), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n523), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n464), .A2(G217), .A3(new_n324), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n535), .B2(new_n544), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n237), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G478), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n550), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n324), .A2(G952), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(G234), .B2(G237), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n324), .B(new_n237), .C1(G234), .C2(G237), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT21), .B(G898), .Z(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n323), .A2(new_n324), .A3(G214), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n514), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(G143), .B2(new_n561), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT18), .A2(G131), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n210), .B(G146), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G113), .B(G122), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n376), .ZN(new_n572));
  INV_X1    g386(.A(new_n223), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n563), .A2(new_n275), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT17), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n563), .B(new_n275), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n573), .B(new_n575), .C1(new_n576), .C2(KEYINPUT17), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n572), .B1(new_n570), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n254), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G475), .ZN(new_n582));
  NAND2_X1  g396(.A1(KEYINPUT94), .A2(KEYINPUT19), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n210), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n210), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n576), .B(new_n214), .C1(G146), .C2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n572), .B1(new_n570), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  NOR4_X1   g403(.A1(new_n589), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT20), .ZN(new_n591));
  INV_X1    g405(.A(new_n588), .ZN(new_n592));
  AOI21_X1  g406(.A(G475), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n593), .B2(new_n254), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n582), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n554), .A2(new_n560), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n365), .A2(new_n463), .A3(new_n513), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n548), .B2(new_n549), .ZN(new_n600));
  INV_X1    g414(.A(new_n549), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(KEYINPUT33), .A3(new_n547), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n600), .A2(new_n602), .A3(G478), .A4(new_n237), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n550), .A2(new_n551), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n594), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n593), .A2(new_n591), .A3(new_n254), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n607), .A2(new_n608), .B1(G475), .B2(new_n581), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n560), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n462), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n459), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n513), .ZN(new_n615));
  INV_X1    g429(.A(new_n252), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n346), .A2(new_n347), .ZN(new_n617));
  OAI21_X1  g431(.A(G472), .B1(new_n617), .B2(new_n236), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n349), .A3(new_n618), .ZN(new_n619));
  NOR4_X1   g433(.A1(new_n612), .A2(new_n614), .A3(new_n615), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT34), .B(G104), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  AOI21_X1  g436(.A(new_n462), .B1(new_n456), .B2(new_n458), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n595), .A2(new_n560), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n623), .A2(new_n554), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n626), .A2(new_n615), .A3(new_n619), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n234), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n228), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n250), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n246), .A2(new_n248), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n618), .A2(new_n349), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n463), .A2(new_n637), .A3(new_n513), .A4(new_n596), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n556), .B1(new_n557), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n553), .A2(new_n595), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n513), .A2(new_n459), .A3(new_n613), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n350), .B(new_n255), .C1(new_n346), .C2(new_n347), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT72), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n350), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n364), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n633), .B(KEYINPUT98), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XOR2_X1   g466(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n642), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n513), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n460), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n609), .A2(new_n553), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n462), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n342), .A2(new_n360), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n329), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n360), .A2(new_n356), .A3(new_n328), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  AOI21_X1  g480(.A(G902), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n663), .B2(new_n664), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n253), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n633), .B1(new_n355), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n656), .A2(new_n658), .A3(new_n661), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n514), .ZN(G45));
  AND3_X1   g487(.A1(new_n513), .A2(new_n613), .A3(new_n459), .ZN(new_n674));
  INV_X1    g488(.A(new_n642), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n605), .A2(new_n595), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n649), .A2(new_n674), .A3(new_n650), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NOR2_X1   g493(.A1(new_n614), .A2(new_n612), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n510), .A2(new_n237), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  INV_X1    g496(.A(new_n465), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n512), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n680), .A2(new_n649), .A3(new_n616), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND3_X1  g502(.A1(new_n365), .A2(new_n625), .A3(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NOR2_X1   g504(.A1(new_n614), .A2(new_n684), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n649), .A3(new_n596), .A4(new_n650), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n635), .B1(new_n364), .B2(new_n355), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(KEYINPUT102), .A3(new_n596), .A4(new_n691), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NOR2_X1   g512(.A1(new_n614), .A2(new_n660), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n339), .B(new_n343), .C1(new_n328), .C2(new_n357), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n253), .A3(new_n254), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n616), .A2(new_n618), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n699), .A2(new_n611), .A3(new_n685), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NAND3_X1  g519(.A1(new_n618), .A2(new_n633), .A3(new_n701), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n691), .A2(new_n677), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  INV_X1    g523(.A(new_n646), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n364), .A2(new_n351), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(KEYINPUT104), .A3(new_n616), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT104), .B1(new_n711), .B2(new_n616), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT42), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n460), .A2(new_n513), .A3(new_n613), .A4(new_n677), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n649), .A2(new_n616), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(new_n716), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT92), .B1(new_n456), .B2(new_n458), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n723), .A2(new_n462), .A3(new_n455), .A4(new_n676), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n365), .A2(new_n513), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(KEYINPUT103), .A3(new_n718), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n717), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n275), .ZN(G33));
  NAND3_X1  g542(.A1(new_n460), .A2(new_n513), .A3(new_n613), .ZN(new_n729));
  INV_X1    g543(.A(new_n643), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n729), .B1(KEYINPUT105), .B2(new_n730), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n365), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  OR2_X1    g548(.A1(new_n503), .A2(new_n487), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(new_n493), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n505), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n512), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT46), .B1(new_n739), .B2(new_n505), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n683), .A4(new_n654), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n609), .A2(new_n605), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n745), .A2(new_n746), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n749), .B2(new_n747), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n636), .A3(new_n633), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(KEYINPUT44), .A3(new_n636), .A4(new_n633), .ZN(new_n756));
  INV_X1    g570(.A(new_n460), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n462), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n683), .B(new_n654), .C1(new_n741), .C2(new_n742), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n744), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  OAI21_X1  g578(.A(new_n683), .B1(new_n741), .B2(new_n742), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(KEYINPUT108), .B2(KEYINPUT47), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n649), .A2(new_n616), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n683), .B(new_n768), .C1(new_n741), .C2(new_n742), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n724), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(new_n658), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n462), .A3(new_n685), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n752), .A2(new_n556), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n703), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT118), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT118), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n773), .A2(new_n775), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n782), .B(new_n776), .C1(new_n773), .C2(new_n775), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n778), .B(new_n779), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n758), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n684), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(new_n707), .A3(new_n774), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n669), .B1(new_n353), .B2(new_n354), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n556), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n616), .A3(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n595), .A3(new_n605), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n786), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n766), .A2(new_n769), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n682), .A2(new_n512), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n683), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n775), .A2(new_n787), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n799), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT116), .A3(new_n465), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT116), .B1(new_n803), .B2(new_n465), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n786), .A2(new_n790), .A3(new_n807), .A4(new_n795), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n796), .A2(new_n802), .B1(new_n808), .B2(new_n797), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n689), .A2(new_n686), .A3(new_n704), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n697), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n727), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n623), .A2(new_n513), .A3(new_n675), .A4(new_n659), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n814), .A2(new_n791), .A3(new_n815), .A4(new_n633), .ZN(new_n816));
  INV_X1    g630(.A(new_n814), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT111), .B1(new_n671), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n678), .A2(new_n651), .A3(new_n708), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n670), .B1(new_n647), .B2(new_n648), .ZN(new_n823));
  INV_X1    g637(.A(new_n633), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n815), .B1(new_n825), .B2(new_n814), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n671), .A2(new_n817), .A3(KEYINPUT111), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n678), .A2(new_n651), .A3(new_n708), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT112), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n822), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n553), .A2(KEYINPUT109), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n553), .A2(KEYINPUT109), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n649), .A2(new_n650), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n595), .A2(new_n642), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n729), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT110), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n836), .A2(new_n729), .A3(new_n842), .A4(new_n839), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n733), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n610), .B1(new_n834), .B2(new_n609), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n845), .A2(new_n615), .A3(new_n619), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n611), .A3(new_n463), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n724), .A2(new_n513), .A3(new_n707), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n597), .A3(new_n638), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT52), .B1(new_n819), .B2(new_n820), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n812), .A2(new_n831), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT112), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT112), .B1(new_n828), .B2(new_n829), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT52), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n812), .A3(new_n831), .A4(new_n850), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n852), .A2(KEYINPUT53), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n857), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n831), .B(new_n851), .C1(new_n812), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n722), .A2(new_n726), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n715), .A2(new_n716), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n810), .A2(new_n697), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n862), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n856), .A2(new_n872), .A3(new_n857), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n861), .A2(new_n870), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n713), .A2(new_n714), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n788), .A2(new_n875), .A3(new_n774), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT48), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n555), .B(KEYINPUT119), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n774), .A2(new_n691), .A3(new_n703), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n788), .A2(new_n616), .A3(new_n610), .A4(new_n792), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT120), .Z(new_n882));
  NAND4_X1  g696(.A1(new_n809), .A2(new_n859), .A3(new_n874), .A4(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n885), .A2(new_n465), .A3(new_n462), .A4(new_n748), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n252), .B1(new_n799), .B2(KEYINPUT49), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n772), .A2(new_n791), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(G75));
  NAND3_X1  g703(.A1(new_n861), .A2(new_n870), .A3(new_n873), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n236), .A3(new_n454), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n450), .B(new_n451), .Z(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n891), .B2(new_n892), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n324), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G51));
  XOR2_X1   g712(.A(new_n505), .B(KEYINPUT57), .Z(new_n899));
  AND3_X1   g713(.A1(new_n856), .A2(new_n872), .A3(new_n857), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n872), .B1(new_n856), .B2(new_n857), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n871), .B1(new_n902), .B2(new_n870), .ZN(new_n903));
  INV_X1    g717(.A(new_n874), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n510), .ZN(new_n906));
  INV_X1    g720(.A(new_n739), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n890), .A2(new_n236), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n897), .B1(new_n906), .B2(new_n908), .ZN(G54));
  NAND4_X1  g723(.A1(new_n890), .A2(KEYINPUT58), .A3(G475), .A4(new_n236), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(new_n589), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n589), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n897), .ZN(G60));
  INV_X1    g727(.A(new_n897), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n874), .B2(new_n859), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n600), .A2(new_n602), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n903), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n921), .B2(new_n874), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(new_n919), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT121), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n890), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n249), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n890), .A2(new_n631), .A3(new_n926), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n914), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n929), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  NAND4_X1  g749(.A1(new_n867), .A2(new_n597), .A3(new_n638), .A4(new_n847), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n324), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT122), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n324), .B1(new_n558), .B2(G224), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n450), .B1(G898), .B2(new_n324), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(G69));
  AND2_X1   g756(.A1(new_n875), .A2(new_n699), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n762), .B(new_n744), .C1(new_n759), .C2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(new_n866), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n770), .A2(new_n733), .A3(new_n829), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n324), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n641), .A2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT124), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n341), .A2(new_n332), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n586), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n672), .A2(new_n829), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n719), .A2(new_n729), .A3(new_n845), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n654), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n960), .A2(new_n763), .A3(new_n770), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n963), .B2(new_n324), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  INV_X1    g779(.A(G227), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n966), .B2(new_n641), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n957), .A2(new_n965), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n955), .B1(new_n950), .B2(new_n952), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n964), .B(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT126), .B(new_n967), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n970), .A2(new_n974), .ZN(G72));
  NOR3_X1   g789(.A1(new_n948), .A2(new_n949), .A3(new_n936), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n361), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n963), .B2(new_n936), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n663), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n361), .A2(new_n979), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n858), .B(new_n985), .C1(new_n662), .C2(new_n329), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n914), .A2(new_n980), .A3(new_n984), .A4(new_n986), .ZN(G57));
endmodule


