//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(G43gat), .A2(G50gat), .ZN(new_n208));
  XOR2_X1   g007(.A(KEYINPUT90), .B(G43gat), .Z(new_n209));
  OAI211_X1 g008(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(G50gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT88), .B(G29gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n211), .A2(G36gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n208), .ZN(new_n217));
  NOR2_X1   g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT15), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n218), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n207), .B1(new_n222), .B2(new_n208), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT89), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n210), .A2(new_n216), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n211), .A2(G36gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n215), .B1(new_n214), .B2(KEYINPUT87), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(new_n212), .B2(new_n213), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n226), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n223), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n206), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(KEYINPUT17), .ZN(new_n234));
  INV_X1    g033(.A(new_n206), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n206), .B(new_n232), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n237), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n237), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT11), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(new_n252), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G22gat), .B(G50gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G228gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n262));
  AND2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264));
  NOR2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G141gat), .B(G148gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G148gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G141gat), .ZN(new_n275));
  INV_X1    g074(.A(G141gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G148gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n265), .A2(KEYINPUT74), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n265), .A2(KEYINPUT74), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n263), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n284));
  NOR2_X1   g083(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n272), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT76), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT76), .B(new_n272), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n278), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n280), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT22), .B1(new_n296), .B2(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n293), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n302));
  INV_X1    g101(.A(G211gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(G218gat), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n292), .A3(new_n298), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n292), .B1(new_n308), .B2(new_n298), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n311), .B2(KEYINPUT79), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n291), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n290), .A2(new_n283), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n266), .A2(new_n262), .A3(new_n267), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT77), .B1(new_n273), .B2(new_n278), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n320), .A3(new_n314), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n261), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT80), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n326), .B(new_n261), .C1(new_n315), .C2(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT31), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT29), .B1(new_n291), .B2(new_n314), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT81), .ZN(new_n331));
  INV_X1    g130(.A(new_n316), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n321), .A2(new_n322), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n314), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n320), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n261), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n328), .A2(new_n329), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n329), .B1(new_n328), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n260), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT65), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n346), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n350), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G190gat), .ZN(new_n353));
  AND2_X1   g152(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT28), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n353), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n352), .A2(new_n357), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G183gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n353), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  INV_X1    g169(.A(G176gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n249), .A2(new_n371), .A3(KEYINPUT23), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(G169gat), .B2(G176gat), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n372), .A2(new_n374), .A3(new_n348), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT64), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n377), .A3(new_n363), .ZN(new_n378));
  OAI211_X1 g177(.A(G183gat), .B(G190gat), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n378), .A2(new_n379), .A3(new_n368), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n374), .A3(new_n348), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT25), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT66), .ZN(new_n385));
  OR2_X1    g184(.A1(G127gat), .A2(G134gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(G127gat), .A2(G134gat), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n384), .A2(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G120gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(G113gat), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT1), .B1(new_n390), .B2(KEYINPUT66), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n389), .A2(G113gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n390), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n386), .A2(new_n387), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n388), .A2(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n344), .B1(new_n383), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT25), .B1(new_n366), .B2(new_n368), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n379), .A3(new_n368), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n375), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n375), .A2(new_n399), .B1(new_n401), .B2(KEYINPUT25), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(KEYINPUT67), .A3(new_n396), .A4(new_n362), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n397), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT68), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT69), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(G71gat), .ZN(new_n412));
  INV_X1    g211(.A(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n407), .A2(new_n417), .A3(KEYINPUT32), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n407), .B(KEYINPUT32), .C1(new_n415), .C2(new_n414), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n405), .A2(new_n406), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT34), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n310), .B2(new_n312), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n330), .A2(new_n316), .B1(new_n427), .B2(new_n291), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n326), .B1(new_n428), .B2(new_n261), .ZN(new_n429));
  INV_X1    g228(.A(new_n327), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n340), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT31), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n328), .A2(new_n329), .A3(new_n340), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n259), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n424), .A2(new_n419), .A3(new_n420), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n343), .A2(new_n426), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  INV_X1    g236(.A(G64gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(G92gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n322), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n383), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n362), .A2(new_n376), .A3(new_n382), .A4(new_n443), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n316), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n316), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n332), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT72), .A3(new_n447), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n440), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n447), .A3(new_n440), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n317), .A2(new_n320), .A3(new_n396), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT4), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n317), .A2(new_n320), .A3(new_n463), .A4(new_n396), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n397), .A3(new_n321), .ZN(new_n467));
  NAND2_X1  g266(.A1(G225gat), .A2(G233gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  INV_X1    g269(.A(new_n461), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n396), .B1(new_n317), .B2(new_n320), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G1gat), .B(G29gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT0), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(G57gat), .ZN(new_n478));
  INV_X1    g277(.A(G85gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT5), .A4(new_n468), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n396), .B1(new_n291), .B2(new_n314), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n487), .A2(new_n466), .B1(new_n462), .B2(new_n464), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n488), .A2(new_n468), .B1(KEYINPUT5), .B2(new_n473), .ZN(new_n489));
  INV_X1    g288(.A(new_n482), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n484), .A3(new_n483), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n436), .A2(new_n460), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  INV_X1    g297(.A(new_n436), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n458), .A2(KEYINPUT73), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT73), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n454), .B2(new_n457), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n502), .A3(new_n459), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n492), .A2(KEYINPUT78), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n491), .A2(new_n505), .A3(new_n484), .A4(new_n483), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n503), .B1(new_n507), .B2(new_n486), .ZN(new_n508));
  AOI211_X1 g307(.A(new_n498), .B(new_n494), .C1(new_n499), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n486), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n341), .A2(new_n342), .A3(new_n260), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n259), .B1(new_n432), .B2(new_n433), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n503), .ZN(new_n514));
  INV_X1    g313(.A(new_n435), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n424), .B1(new_n420), .B2(new_n419), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n510), .A2(new_n513), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT86), .B1(new_n518), .B2(KEYINPUT35), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n497), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n465), .A2(new_n467), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT82), .B(KEYINPUT39), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n470), .A3(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n471), .A2(new_n472), .A3(new_n470), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT83), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n488), .B2(new_n468), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT39), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n480), .B(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT40), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT40), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(KEYINPUT84), .A3(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n531), .A2(new_n483), .A3(new_n533), .A4(new_n460), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n450), .B2(new_n453), .ZN(new_n537));
  INV_X1    g336(.A(new_n440), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n452), .A2(new_n447), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(KEYINPUT37), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT38), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n537), .C2(new_n540), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n455), .A3(new_n544), .ZN(new_n545));
  AOI211_X1 g344(.A(KEYINPUT38), .B(new_n540), .C1(new_n539), .C2(KEYINPUT37), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n545), .A2(new_n546), .A3(new_n493), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n535), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n510), .A2(new_n514), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n343), .A2(new_n434), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n515), .B2(new_n516), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n426), .A2(KEYINPUT36), .A3(new_n435), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n256), .B1(new_n520), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G57gat), .ZN(new_n558));
  OR3_X1    g357(.A1(new_n558), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(new_n558), .B2(G64gat), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n559), .B(new_n560), .C1(G57gat), .C2(new_n438), .ZN(new_n561));
  NAND2_X1  g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  OR2_X1    g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n562), .B(KEYINPUT91), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n564), .A2(KEYINPUT91), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n567), .B(new_n563), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n206), .B1(KEYINPUT21), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT19), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT93), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n571), .A2(KEYINPUT21), .ZN(new_n578));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n578), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n577), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n479), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT94), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT7), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(new_n592), .C1(new_n587), .C2(new_n586), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT96), .B(G92gat), .Z(new_n594));
  INV_X1    g393(.A(KEYINPUT8), .ZN(new_n595));
  NOR2_X1   g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n594), .A2(new_n479), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n593), .B(new_n600), .C1(new_n592), .C2(new_n591), .ZN(new_n601));
  INV_X1    g400(.A(new_n596), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT97), .B1(new_n602), .B2(new_n599), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(new_n571), .Z(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n571), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n605), .A2(new_n610), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n371), .ZN(new_n615));
  INV_X1    g414(.A(G204gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n613), .B2(new_n618), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n232), .ZN(new_n625));
  NAND3_X1  g424(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n232), .B(KEYINPUT17), .Z(new_n627));
  OAI211_X1 g426(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n604), .ZN(new_n628));
  XOR2_X1   g427(.A(G190gat), .B(G218gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT98), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n634), .B1(new_n633), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n639), .A2(new_n631), .A3(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n584), .A2(new_n624), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n557), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n485), .B1(new_n504), .B2(new_n506), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n460), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  MUX2_X1   g454(.A(new_n653), .B(new_n655), .S(KEYINPUT42), .Z(G1325gat));
  XNOR2_X1  g455(.A(new_n555), .B(KEYINPUT101), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n646), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n426), .A2(new_n435), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT102), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n513), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n644), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n520), .B2(new_n556), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n624), .A2(new_n583), .A3(new_n256), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n669), .A2(new_n510), .A3(new_n211), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT45), .Z(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n436), .A2(new_n648), .A3(new_n503), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n498), .B1(new_n674), .B2(new_n494), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n518), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n496), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n549), .B2(new_n550), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n555), .B1(new_n535), .B2(new_n547), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n678), .B(new_n550), .C1(new_n648), .C2(new_n503), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n673), .B(new_n644), .C1(new_n677), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n667), .B2(new_n673), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(new_n668), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n672), .B1(new_n687), .B2(new_n510), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(KEYINPUT104), .A3(new_n648), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n211), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n671), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT105), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n694), .B(new_n671), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1328gat));
  INV_X1    g495(.A(new_n460), .ZN(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n687), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n669), .A2(G36gat), .A3(new_n697), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(new_n209), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n667), .A2(new_n703), .A3(new_n517), .A4(new_n668), .ZN(new_n704));
  INV_X1    g503(.A(new_n555), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n686), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT108), .ZN(new_n707));
  OAI211_X1 g506(.A(KEYINPUT47), .B(new_n704), .C1(new_n707), .C2(new_n703), .ZN(new_n708));
  INV_X1    g507(.A(new_n657), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n703), .B1(new_n686), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n704), .B(KEYINPUT107), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(KEYINPUT47), .B2(new_n712), .ZN(G1330gat));
  OAI21_X1  g512(.A(G50gat), .B1(new_n687), .B2(new_n513), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT48), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n669), .B(KEYINPUT109), .ZN(new_n717));
  INV_X1    g516(.A(G50gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n550), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n716), .B(new_n720), .ZN(G1331gat));
  NAND2_X1  g520(.A1(new_n551), .A2(KEYINPUT103), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n722), .A2(new_n548), .A3(new_n555), .A4(new_n681), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n584), .B1(new_n520), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n613), .A2(new_n618), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n622), .B2(new_n619), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n256), .B1(new_n642), .B2(new_n643), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n510), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n558), .ZN(G1332gat));
  INV_X1    g530(.A(new_n729), .ZN(new_n732));
  NAND2_X1  g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n460), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT111), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n732), .B2(new_n709), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n729), .A2(new_n659), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT112), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n739), .B1(new_n741), .B2(new_n738), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n550), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n583), .A2(new_n255), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n624), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT113), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n685), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n749), .A2(new_n479), .A3(new_n510), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n644), .B(new_n746), .C1(new_n677), .C2(new_n683), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n520), .A2(new_n723), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n644), .A4(new_n746), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n726), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n648), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n750), .A2(new_n757), .ZN(G1336gat));
  INV_X1    g557(.A(new_n594), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n749), .B2(new_n697), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n585), .A3(new_n460), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n749), .B2(new_n657), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n753), .A2(new_n755), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n624), .A2(new_n413), .A3(new_n517), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT115), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n685), .A2(new_n550), .A3(new_n748), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n513), .A2(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT116), .B1(new_n776), .B2(KEYINPUT53), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n778), .B(new_n779), .C1(new_n773), .C2(new_n775), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781));
  AOI22_X1  g580(.A1(G106gat), .A2(new_n772), .B1(new_n756), .B2(new_n774), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n783));
  AOI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND4_X1   g583(.A1(new_n781), .A2(new_n773), .A3(new_n775), .A4(new_n783), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n777), .A2(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n778), .B1(new_n782), .B2(new_n779), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n776), .A2(KEYINPUT116), .A3(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(KEYINPUT119), .C1(new_n784), .C2(new_n785), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1339gat));
  NOR2_X1   g592(.A1(new_n236), .A2(new_n237), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n241), .A2(new_n242), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n250), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n253), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n644), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n617), .B1(new_n611), .B2(KEYINPUT54), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n607), .A2(G230gat), .A3(G233gat), .A4(new_n608), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n611), .A2(KEYINPUT54), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n803), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT55), .B1(new_n805), .B2(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n798), .A2(new_n623), .A3(new_n807), .A4(new_n727), .ZN(new_n808));
  INV_X1    g607(.A(new_n797), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n624), .A2(new_n666), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n583), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n583), .A2(new_n666), .A3(new_n726), .A4(new_n256), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n648), .B(new_n697), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n436), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n255), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n624), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n583), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(G127gat), .ZN(G1342gat));
  NOR3_X1   g619(.A1(new_n813), .A2(new_n666), .A3(new_n436), .ZN(new_n821));
  NOR2_X1   g620(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n822));
  AND2_X1   g621(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n821), .B2(new_n822), .ZN(G1343gat));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n810), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n812), .B1(new_n827), .B2(new_n584), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(new_n513), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT57), .B(new_n550), .C1(new_n811), .C2(new_n812), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n705), .A2(new_n510), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n697), .A3(new_n255), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G141gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n657), .A2(new_n550), .ZN(new_n835));
  NOR4_X1   g634(.A1(new_n813), .A2(G141gat), .A3(new_n835), .A4(new_n256), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT58), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n834), .B2(new_n837), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT120), .B(new_n836), .C1(new_n833), .C2(G141gat), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n842), .A2(new_n846), .ZN(G1344gat));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n697), .A3(new_n832), .ZN(new_n848));
  OAI21_X1  g647(.A(G148gat), .B1(new_n848), .B2(new_n726), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n813), .A2(new_n835), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n274), .A3(new_n624), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT121), .Z(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(G1345gat));
  OAI21_X1  g655(.A(G155gat), .B1(new_n848), .B2(new_n584), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n269), .A3(new_n583), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1346gat));
  OAI21_X1  g658(.A(G162gat), .B1(new_n848), .B2(new_n666), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n853), .A2(new_n270), .A3(new_n644), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1347gat));
  NOR3_X1   g661(.A1(new_n828), .A2(new_n648), .A3(new_n697), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n499), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n256), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(new_n249), .ZN(G1348gat));
  NAND2_X1  g665(.A1(KEYINPUT122), .A2(G176gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(new_n864), .B2(new_n726), .ZN(new_n868));
  NOR2_X1   g667(.A1(KEYINPUT122), .A2(G176gat), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1349gat));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT123), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n367), .B1(new_n864), .B2(new_n584), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n863), .A2(new_n583), .A3(new_n499), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n359), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n871), .A2(KEYINPUT123), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n875), .B(new_n876), .Z(G1350gat));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G190gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n666), .ZN(new_n880));
  MUX2_X1   g679(.A(new_n878), .B(new_n879), .S(new_n880), .Z(G1351gat));
  NAND4_X1  g680(.A1(new_n831), .A2(new_n510), .A3(new_n460), .A4(new_n657), .ZN(new_n882));
  OAI21_X1  g681(.A(G197gat), .B1(new_n882), .B2(new_n256), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n550), .A3(new_n657), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n256), .A2(G197gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1352gat));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n884), .A2(G204gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n624), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n884), .A2(KEYINPUT124), .A3(G204gat), .A4(new_n726), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n882), .A2(KEYINPUT125), .A3(new_n726), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT125), .B1(new_n882), .B2(new_n726), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(G204gat), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(G1353gat));
  OR2_X1    g696(.A1(new_n882), .A2(new_n584), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G211gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT63), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n884), .A2(new_n584), .A3(new_n296), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n900), .A2(KEYINPUT63), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(KEYINPUT63), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n898), .A2(G211gat), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(G1354gat));
  OR2_X1    g705(.A1(new_n882), .A2(KEYINPUT127), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n882), .A2(KEYINPUT127), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n644), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G218gat), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n666), .A2(G218gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n884), .B2(new_n911), .ZN(G1355gat));
endmodule


