

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734;

  INV_X1 U374 ( .A(G146), .ZN(n362) );
  XNOR2_X1 U375 ( .A(n533), .B(KEYINPUT45), .ZN(n705) );
  NOR2_X1 U376 ( .A1(n562), .A2(n653), .ZN(n564) );
  INV_X1 U377 ( .A(n580), .ZN(n375) );
  XNOR2_X2 U378 ( .A(n510), .B(KEYINPUT1), .ZN(n575) );
  OR2_X1 U379 ( .A1(n645), .A2(n552), .ZN(n560) );
  BUF_X1 U380 ( .A(n490), .Z(n442) );
  INV_X2 U381 ( .A(G953), .ZN(n704) );
  XNOR2_X2 U382 ( .A(G119), .B(G110), .ZN(n355) );
  XNOR2_X2 U383 ( .A(n384), .B(KEYINPUT0), .ZN(n514) );
  XOR2_X2 U384 ( .A(KEYINPUT10), .B(n387), .Z(n427) );
  XNOR2_X2 U385 ( .A(n362), .B(G125), .ZN(n387) );
  INV_X1 U386 ( .A(G110), .ZN(n417) );
  NAND2_X1 U387 ( .A1(n502), .A2(n353), .ZN(n509) );
  AND2_X2 U388 ( .A1(n597), .A2(n596), .ZN(n689) );
  INV_X1 U389 ( .A(n595), .ZN(n596) );
  XNOR2_X1 U390 ( .A(n418), .B(n417), .ZN(n419) );
  AND2_X1 U391 ( .A1(n603), .A2(G953), .ZN(n703) );
  AND2_X1 U392 ( .A1(n501), .A2(n528), .ZN(n353) );
  XNOR2_X2 U393 ( .A(n425), .B(n424), .ZN(n510) );
  XOR2_X1 U394 ( .A(KEYINPUT78), .B(KEYINPUT8), .Z(n354) );
  NAND2_X1 U395 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U396 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U397 ( .A(G143), .B(G128), .ZN(n406) );
  NOR2_X1 U398 ( .A1(n637), .A2(n537), .ZN(n576) );
  AND2_X1 U399 ( .A1(n587), .A2(n586), .ZN(n724) );
  XNOR2_X1 U400 ( .A(n420), .B(n419), .ZN(n423) );
  OR2_X1 U401 ( .A1(n653), .A2(n464), .ZN(n466) );
  XNOR2_X1 U402 ( .A(n401), .B(n400), .ZN(n517) );
  XOR2_X1 U403 ( .A(n517), .B(KEYINPUT97), .Z(n522) );
  OR2_X1 U404 ( .A1(n486), .A2(n575), .ZN(n462) );
  XOR2_X1 U405 ( .A(G116), .B(G107), .Z(n409) );
  XNOR2_X1 U406 ( .A(KEYINPUT16), .B(n355), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n409), .B(n356), .ZN(n358) );
  XNOR2_X1 U408 ( .A(G113), .B(G104), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n357), .B(G122), .ZN(n388) );
  XNOR2_X1 U410 ( .A(n358), .B(n388), .ZN(n710) );
  NAND2_X1 U411 ( .A1(n704), .A2(G224), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n359), .B(KEYINPUT73), .ZN(n361) );
  XNOR2_X1 U413 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n363), .B(n387), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n710), .B(n364), .ZN(n368) );
  XNOR2_X1 U417 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n406), .B(n365), .ZN(n722) );
  INV_X1 U419 ( .A(G101), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n722), .B(n366), .ZN(n421) );
  INV_X1 U421 ( .A(KEYINPUT67), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n367), .B(KEYINPUT3), .ZN(n712) );
  XNOR2_X1 U423 ( .A(n421), .B(n712), .ZN(n454) );
  XNOR2_X1 U424 ( .A(n368), .B(n454), .ZN(n609) );
  XNOR2_X1 U425 ( .A(KEYINPUT15), .B(G902), .ZN(n595) );
  NAND2_X1 U426 ( .A1(n609), .A2(n595), .ZN(n373) );
  INV_X1 U427 ( .A(G902), .ZN(n456) );
  INV_X1 U428 ( .A(G237), .ZN(n369) );
  NAND2_X1 U429 ( .A1(n456), .A2(n369), .ZN(n374) );
  NAND2_X1 U430 ( .A1(n374), .A2(G210), .ZN(n371) );
  INV_X1 U431 ( .A(KEYINPUT85), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X2 U433 ( .A(n373), .B(n372), .ZN(n580) );
  NAND2_X1 U434 ( .A1(n374), .A2(G214), .ZN(n649) );
  INV_X1 U435 ( .A(n649), .ZN(n652) );
  NAND2_X1 U436 ( .A1(n375), .A2(n649), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n376), .B(KEYINPUT19), .ZN(n554) );
  NAND2_X1 U438 ( .A1(G234), .A2(G237), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n377), .B(KEYINPUT86), .ZN(n378) );
  XNOR2_X1 U440 ( .A(KEYINPUT14), .B(n378), .ZN(n380) );
  NAND2_X1 U441 ( .A1(n380), .A2(G902), .ZN(n379) );
  XOR2_X1 U442 ( .A(KEYINPUT88), .B(n379), .Z(n468) );
  NOR2_X1 U443 ( .A1(G898), .A2(n704), .ZN(n715) );
  NAND2_X1 U444 ( .A1(n468), .A2(n715), .ZN(n382) );
  NAND2_X1 U445 ( .A1(n380), .A2(G952), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n381), .B(KEYINPUT87), .ZN(n678) );
  NAND2_X1 U447 ( .A1(n678), .A2(n704), .ZN(n467) );
  NAND2_X1 U448 ( .A1(n382), .A2(n467), .ZN(n383) );
  NAND2_X1 U449 ( .A1(n554), .A2(n383), .ZN(n384) );
  NAND2_X1 U450 ( .A1(G234), .A2(n595), .ZN(n385) );
  XNOR2_X1 U451 ( .A(KEYINPUT20), .B(n385), .ZN(n438) );
  AND2_X1 U452 ( .A1(n438), .A2(G221), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n386), .B(KEYINPUT21), .ZN(n663) );
  XNOR2_X1 U454 ( .A(KEYINPUT13), .B(G475), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n388), .B(n427), .ZN(n389) );
  INV_X1 U456 ( .A(n389), .ZN(n391) );
  NOR2_X1 U457 ( .A1(G953), .A2(G237), .ZN(n449) );
  NAND2_X1 U458 ( .A1(G214), .A2(n449), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n399) );
  XOR2_X1 U460 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n393) );
  XNOR2_X1 U461 ( .A(G143), .B(KEYINPUT94), .ZN(n392) );
  XNOR2_X1 U462 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U463 ( .A(G140), .B(KEYINPUT96), .Z(n395) );
  XNOR2_X1 U464 ( .A(G131), .B(KEYINPUT11), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U466 ( .A(n397), .B(n396), .Z(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n600) );
  NOR2_X1 U468 ( .A1(G902), .A2(n600), .ZN(n400) );
  XOR2_X1 U469 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n404) );
  NAND2_X1 U470 ( .A1(G234), .A2(n704), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n354), .B(n402), .ZN(n434) );
  NAND2_X1 U472 ( .A1(G217), .A2(n434), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U474 ( .A(G122), .B(G134), .Z(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U476 ( .A(n408), .B(n407), .Z(n411) );
  XNOR2_X1 U477 ( .A(n409), .B(KEYINPUT9), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n697) );
  NOR2_X1 U479 ( .A1(G902), .A2(n697), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n412), .B(G478), .ZN(n521) );
  INV_X1 U481 ( .A(n521), .ZN(n518) );
  NOR2_X1 U482 ( .A1(n517), .A2(n518), .ZN(n654) );
  NAND2_X1 U483 ( .A1(n663), .A2(n654), .ZN(n413) );
  OR2_X2 U484 ( .A1(n514), .A2(n413), .ZN(n414) );
  XNOR2_X1 U485 ( .A(n414), .B(KEYINPUT22), .ZN(n486) );
  XNOR2_X1 U486 ( .A(G137), .B(G140), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n426), .B(G107), .ZN(n416) );
  XNOR2_X1 U488 ( .A(G131), .B(G134), .ZN(n721) );
  XNOR2_X1 U489 ( .A(n721), .B(G146), .ZN(n443) );
  XNOR2_X1 U490 ( .A(n443), .B(G104), .ZN(n415) );
  XNOR2_X1 U491 ( .A(n416), .B(n415), .ZN(n420) );
  NAND2_X1 U492 ( .A1(G227), .A2(n704), .ZN(n418) );
  INV_X1 U493 ( .A(n421), .ZN(n422) );
  XNOR2_X1 U494 ( .A(n423), .B(n422), .ZN(n693) );
  NAND2_X1 U495 ( .A1(n693), .A2(n456), .ZN(n425) );
  XNOR2_X1 U496 ( .A(KEYINPUT66), .B(G469), .ZN(n424) );
  XNOR2_X1 U497 ( .A(n462), .B(KEYINPUT103), .ZN(n459) );
  XNOR2_X1 U498 ( .A(n427), .B(n426), .ZN(n719) );
  XOR2_X1 U499 ( .A(G119), .B(G110), .Z(n428) );
  XNOR2_X1 U500 ( .A(G128), .B(n428), .ZN(n429) );
  XNOR2_X1 U501 ( .A(n429), .B(KEYINPUT24), .ZN(n433) );
  XOR2_X1 U502 ( .A(KEYINPUT72), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U503 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n430) );
  XNOR2_X1 U504 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U505 ( .A(n433), .B(n432), .Z(n436) );
  NAND2_X1 U506 ( .A1(G221), .A2(n434), .ZN(n435) );
  XNOR2_X1 U507 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U508 ( .A(n719), .B(n437), .ZN(n700) );
  NOR2_X1 U509 ( .A1(n700), .A2(G902), .ZN(n441) );
  NAND2_X1 U510 ( .A1(n438), .A2(G217), .ZN(n439) );
  XNOR2_X1 U511 ( .A(KEYINPUT25), .B(n439), .ZN(n440) );
  XNOR2_X1 U512 ( .A(n441), .B(n440), .ZN(n490) );
  XOR2_X1 U513 ( .A(KEYINPUT70), .B(G113), .Z(n445) );
  XNOR2_X1 U514 ( .A(G119), .B(G116), .ZN(n444) );
  XNOR2_X1 U515 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U516 ( .A(n443), .B(n446), .ZN(n453) );
  XOR2_X1 U517 ( .A(G137), .B(KEYINPUT91), .Z(n448) );
  XNOR2_X1 U518 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n447) );
  XNOR2_X1 U519 ( .A(n448), .B(n447), .ZN(n451) );
  NAND2_X1 U520 ( .A1(n449), .A2(G210), .ZN(n450) );
  XNOR2_X1 U521 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U522 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U523 ( .A(n455), .B(n454), .ZN(n614) );
  NAND2_X1 U524 ( .A1(n614), .A2(n456), .ZN(n457) );
  XNOR2_X2 U525 ( .A(n457), .B(G472), .ZN(n542) );
  NOR2_X1 U526 ( .A1(n442), .A2(n542), .ZN(n458) );
  NAND2_X1 U527 ( .A1(n459), .A2(n458), .ZN(n503) );
  XNOR2_X1 U528 ( .A(n503), .B(G110), .ZN(G12) );
  XNOR2_X1 U529 ( .A(KEYINPUT6), .B(KEYINPUT100), .ZN(n460) );
  XNOR2_X1 U530 ( .A(n542), .B(n460), .ZN(n535) );
  NAND2_X1 U531 ( .A1(n535), .A2(n442), .ZN(n461) );
  OR2_X1 U532 ( .A1(n462), .A2(n461), .ZN(n524) );
  XNOR2_X1 U533 ( .A(n524), .B(G101), .ZN(G3) );
  XNOR2_X1 U534 ( .A(KEYINPUT69), .B(KEYINPUT38), .ZN(n463) );
  XNOR2_X1 U535 ( .A(n580), .B(n463), .ZN(n653) );
  NAND2_X1 U536 ( .A1(n654), .A2(n649), .ZN(n464) );
  XNOR2_X1 U537 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n465) );
  XNOR2_X1 U538 ( .A(n466), .B(n465), .ZN(n682) );
  INV_X1 U539 ( .A(n467), .ZN(n471) );
  NAND2_X1 U540 ( .A1(G953), .A2(n468), .ZN(n469) );
  NOR2_X1 U541 ( .A1(G900), .A2(n469), .ZN(n470) );
  NOR2_X1 U542 ( .A1(n471), .A2(n470), .ZN(n545) );
  NOR2_X1 U543 ( .A1(n545), .A2(n490), .ZN(n472) );
  NAND2_X1 U544 ( .A1(n472), .A2(n663), .ZN(n534) );
  INV_X1 U545 ( .A(n542), .ZN(n665) );
  NOR2_X1 U546 ( .A1(n534), .A2(n665), .ZN(n475) );
  XNOR2_X1 U547 ( .A(KEYINPUT28), .B(KEYINPUT107), .ZN(n473) );
  XOR2_X1 U548 ( .A(n473), .B(KEYINPUT108), .Z(n474) );
  XNOR2_X1 U549 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U550 ( .A1(n476), .A2(n510), .ZN(n553) );
  OR2_X1 U551 ( .A1(n682), .A2(n553), .ZN(n478) );
  INV_X1 U552 ( .A(KEYINPUT42), .ZN(n477) );
  XNOR2_X1 U553 ( .A(n478), .B(n477), .ZN(n561) );
  XOR2_X1 U554 ( .A(G137), .B(KEYINPUT126), .Z(n479) );
  XNOR2_X1 U555 ( .A(n561), .B(n479), .ZN(G39) );
  INV_X1 U556 ( .A(KEYINPUT82), .ZN(n480) );
  XNOR2_X1 U557 ( .A(n480), .B(n575), .ZN(n541) );
  NOR2_X1 U558 ( .A1(n541), .A2(n442), .ZN(n481) );
  XNOR2_X1 U559 ( .A(KEYINPUT102), .B(n481), .ZN(n483) );
  XNOR2_X1 U560 ( .A(n535), .B(KEYINPUT76), .ZN(n482) );
  AND2_X1 U561 ( .A1(n483), .A2(n482), .ZN(n485) );
  INV_X1 U562 ( .A(KEYINPUT75), .ZN(n484) );
  XNOR2_X1 U563 ( .A(n485), .B(n484), .ZN(n488) );
  INV_X1 U564 ( .A(n486), .ZN(n487) );
  NAND2_X1 U565 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U566 ( .A(n489), .B(KEYINPUT32), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(G119), .ZN(G21) );
  NAND2_X1 U568 ( .A1(n503), .A2(n504), .ZN(n502) );
  NAND2_X1 U569 ( .A1(n663), .A2(n490), .ZN(n660) );
  INV_X1 U570 ( .A(n660), .ZN(n491) );
  NAND2_X1 U571 ( .A1(n575), .A2(n491), .ZN(n513) );
  OR2_X1 U572 ( .A1(n513), .A2(n535), .ZN(n492) );
  XNOR2_X2 U573 ( .A(n492), .B(KEYINPUT33), .ZN(n684) );
  INV_X1 U574 ( .A(n514), .ZN(n493) );
  NAND2_X1 U575 ( .A1(n684), .A2(n493), .ZN(n495) );
  INV_X1 U576 ( .A(KEYINPUT34), .ZN(n494) );
  XNOR2_X1 U577 ( .A(n495), .B(n494), .ZN(n497) );
  NAND2_X1 U578 ( .A1(n517), .A2(n518), .ZN(n548) );
  INV_X1 U579 ( .A(n548), .ZN(n496) );
  NAND2_X1 U580 ( .A1(n497), .A2(n496), .ZN(n500) );
  XNOR2_X1 U581 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n498) );
  XNOR2_X1 U582 ( .A(n498), .B(KEYINPUT74), .ZN(n499) );
  XNOR2_X2 U583 ( .A(n500), .B(n499), .ZN(n621) );
  NAND2_X1 U584 ( .A1(n621), .A2(KEYINPUT81), .ZN(n501) );
  INV_X1 U585 ( .A(KEYINPUT44), .ZN(n528) );
  AND2_X1 U586 ( .A1(n504), .A2(n503), .ZN(n507) );
  NOR2_X1 U587 ( .A1(KEYINPUT81), .A2(KEYINPUT44), .ZN(n505) );
  NAND2_X1 U588 ( .A1(n621), .A2(n505), .ZN(n506) );
  NAND2_X1 U589 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U590 ( .A1(n509), .A2(n508), .ZN(n532) );
  INV_X1 U591 ( .A(KEYINPUT101), .ZN(n527) );
  INV_X1 U592 ( .A(n510), .ZN(n511) );
  NOR2_X1 U593 ( .A1(n511), .A2(n660), .ZN(n547) );
  NAND2_X1 U594 ( .A1(n547), .A2(n665), .ZN(n512) );
  OR2_X1 U595 ( .A1(n514), .A2(n512), .ZN(n623) );
  OR2_X1 U596 ( .A1(n513), .A2(n665), .ZN(n670) );
  NOR2_X1 U597 ( .A1(n514), .A2(n670), .ZN(n516) );
  XOR2_X1 U598 ( .A(KEYINPUT93), .B(KEYINPUT31), .Z(n515) );
  XNOR2_X1 U599 ( .A(n516), .B(n515), .ZN(n639) );
  NAND2_X1 U600 ( .A1(n623), .A2(n639), .ZN(n523) );
  INV_X1 U601 ( .A(n522), .ZN(n519) );
  NAND2_X1 U602 ( .A1(n519), .A2(n518), .ZN(n640) );
  INV_X1 U603 ( .A(KEYINPUT99), .ZN(n520) );
  XNOR2_X1 U604 ( .A(n640), .B(n520), .ZN(n584) );
  NAND2_X1 U605 ( .A1(n522), .A2(n521), .ZN(n637) );
  NAND2_X1 U606 ( .A1(n584), .A2(n637), .ZN(n650) );
  NAND2_X1 U607 ( .A1(n523), .A2(n650), .ZN(n525) );
  NAND2_X1 U608 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U609 ( .A(n527), .B(n526), .ZN(n530) );
  NOR2_X1 U610 ( .A1(n621), .A2(n528), .ZN(n529) );
  NOR2_X1 U611 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U612 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U613 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U614 ( .A1(n536), .A2(n649), .ZN(n537) );
  NAND2_X1 U615 ( .A1(n576), .A2(n375), .ZN(n538) );
  XNOR2_X1 U616 ( .A(n538), .B(KEYINPUT36), .ZN(n539) );
  XNOR2_X1 U617 ( .A(n539), .B(KEYINPUT110), .ZN(n540) );
  NOR2_X1 U618 ( .A1(n541), .A2(n540), .ZN(n645) );
  NAND2_X1 U619 ( .A1(n542), .A2(n649), .ZN(n543) );
  XNOR2_X1 U620 ( .A(KEYINPUT30), .B(n543), .ZN(n544) );
  NOR2_X1 U621 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U622 ( .A1(n547), .A2(n546), .ZN(n562) );
  NOR2_X1 U623 ( .A1(n562), .A2(n548), .ZN(n549) );
  AND2_X1 U624 ( .A1(n549), .A2(n375), .ZN(n633) );
  INV_X1 U625 ( .A(n633), .ZN(n551) );
  INV_X1 U626 ( .A(KEYINPUT68), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n556), .A2(KEYINPUT47), .ZN(n550) );
  NAND2_X1 U628 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U629 ( .A(n553), .ZN(n555) );
  AND2_X1 U630 ( .A1(n555), .A2(n554), .ZN(n635) );
  NAND2_X1 U631 ( .A1(n650), .A2(n635), .ZN(n558) );
  OR2_X1 U632 ( .A1(n556), .A2(KEYINPUT47), .ZN(n557) );
  XNOR2_X1 U633 ( .A(n558), .B(n557), .ZN(n559) );
  NOR2_X1 U634 ( .A1(n560), .A2(n559), .ZN(n572) );
  INV_X1 U635 ( .A(n561), .ZN(n568) );
  XNOR2_X1 U636 ( .A(KEYINPUT80), .B(KEYINPUT39), .ZN(n563) );
  XNOR2_X1 U637 ( .A(n564), .B(n563), .ZN(n585) );
  OR2_X1 U638 ( .A1(n585), .A2(n637), .ZN(n566) );
  INV_X1 U639 ( .A(KEYINPUT40), .ZN(n565) );
  XNOR2_X1 U640 ( .A(n566), .B(n565), .ZN(n732) );
  INV_X1 U641 ( .A(n732), .ZN(n567) );
  INV_X1 U642 ( .A(KEYINPUT46), .ZN(n569) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U644 ( .A(KEYINPUT48), .ZN(n573) );
  XNOR2_X1 U645 ( .A(n574), .B(n573), .ZN(n587) );
  INV_X1 U646 ( .A(n575), .ZN(n661) );
  NAND2_X1 U647 ( .A1(n576), .A2(n661), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n577) );
  XNOR2_X1 U649 ( .A(KEYINPUT105), .B(n577), .ZN(n578) );
  XNOR2_X1 U650 ( .A(n579), .B(n578), .ZN(n581) );
  AND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U652 ( .A(KEYINPUT106), .ZN(n582) );
  XNOR2_X1 U653 ( .A(n583), .B(n582), .ZN(n734) );
  OR2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n646) );
  AND2_X1 U655 ( .A1(n734), .A2(n646), .ZN(n586) );
  NOR2_X1 U656 ( .A1(KEYINPUT2), .A2(KEYINPUT71), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n724), .A2(n588), .ZN(n591) );
  INV_X1 U658 ( .A(n724), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n589), .A2(KEYINPUT71), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n705), .A2(n592), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n705), .A2(n724), .ZN(n648) );
  NAND2_X1 U663 ( .A1(n648), .A2(KEYINPUT2), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n689), .A2(G475), .ZN(n602) );
  XNOR2_X1 U666 ( .A(KEYINPUT83), .B(KEYINPUT121), .ZN(n598) );
  XOR2_X1 U667 ( .A(n598), .B(KEYINPUT59), .Z(n599) );
  XNOR2_X1 U668 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U669 ( .A(n602), .B(n601), .ZN(n604) );
  INV_X1 U670 ( .A(G952), .ZN(n603) );
  NOR2_X2 U671 ( .A1(n604), .A2(n703), .ZN(n606) );
  XNOR2_X1 U672 ( .A(KEYINPUT64), .B(KEYINPUT60), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n606), .B(n605), .ZN(G60) );
  NAND2_X1 U674 ( .A1(n689), .A2(G210), .ZN(n611) );
  XNOR2_X1 U675 ( .A(KEYINPUT77), .B(KEYINPUT54), .ZN(n607) );
  XOR2_X1 U676 ( .A(n607), .B(KEYINPUT55), .Z(n608) );
  XNOR2_X1 U677 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X2 U679 ( .A1(n612), .A2(n703), .ZN(n613) );
  XNOR2_X1 U680 ( .A(n613), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U681 ( .A1(n689), .A2(G472), .ZN(n616) );
  XOR2_X1 U682 ( .A(KEYINPUT62), .B(n614), .Z(n615) );
  XNOR2_X1 U683 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X2 U684 ( .A1(n617), .A2(n703), .ZN(n620) );
  XNOR2_X1 U685 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n618), .B(KEYINPUT84), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(G57) );
  XNOR2_X1 U688 ( .A(n621), .B(G122), .ZN(G24) );
  NOR2_X1 U689 ( .A1(n637), .A2(n623), .ZN(n622) );
  XOR2_X1 U690 ( .A(G104), .B(n622), .Z(G6) );
  NOR2_X1 U691 ( .A1(n640), .A2(n623), .ZN(n628) );
  XOR2_X1 U692 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n625) );
  XNOR2_X1 U693 ( .A(G107), .B(KEYINPUT112), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(KEYINPUT26), .B(n626), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(G9) );
  XOR2_X1 U697 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n631) );
  INV_X1 U698 ( .A(n640), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n635), .A2(n629), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U701 ( .A(G128), .B(n632), .ZN(G30) );
  XOR2_X1 U702 ( .A(G143), .B(n633), .Z(G45) );
  INV_X1 U703 ( .A(n637), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U705 ( .A(G146), .B(n636), .ZN(G48) );
  NOR2_X1 U706 ( .A1(n637), .A2(n639), .ZN(n638) );
  XOR2_X1 U707 ( .A(G113), .B(n638), .Z(G15) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U709 ( .A(G116), .B(n641), .Z(G18) );
  XOR2_X1 U710 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n643) );
  XNOR2_X1 U711 ( .A(G125), .B(KEYINPUT37), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n645), .B(n644), .ZN(G27) );
  INV_X1 U714 ( .A(n646), .ZN(n647) );
  XOR2_X1 U715 ( .A(G134), .B(n647), .Z(G36) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n648), .Z(n681) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n651), .A2(n653), .ZN(n657) );
  NAND2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n655) );
  AND2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n659) );
  INV_X1 U722 ( .A(n684), .ZN(n658) );
  NOR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n676) );
  XNOR2_X1 U724 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n673) );
  NAND2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U726 ( .A(n662), .B(KEYINPUT50), .ZN(n669) );
  NOR2_X1 U727 ( .A1(n663), .A2(n442), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n664), .B(KEYINPUT49), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U730 ( .A(KEYINPUT117), .B(n667), .ZN(n668) );
  NAND2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U733 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U734 ( .A1(n674), .A2(n682), .ZN(n675) );
  NOR2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U736 ( .A(KEYINPUT52), .B(n677), .Z(n679) );
  NAND2_X1 U737 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U738 ( .A1(n681), .A2(n680), .ZN(n687) );
  INV_X1 U739 ( .A(n682), .ZN(n683) );
  NAND2_X1 U740 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U741 ( .A1(n685), .A2(n704), .ZN(n686) );
  NOR2_X1 U742 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U743 ( .A(n688), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U744 ( .A1(n689), .A2(G469), .ZN(n695) );
  XOR2_X1 U745 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n691) );
  XNOR2_X1 U746 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U749 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n703), .A2(n696), .ZN(G54) );
  NAND2_X1 U751 ( .A1(n689), .A2(G478), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U753 ( .A1(n703), .A2(n699), .ZN(G63) );
  NAND2_X1 U754 ( .A1(n689), .A2(G217), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n703), .A2(n702), .ZN(G66) );
  NAND2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U759 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U760 ( .A1(n707), .A2(G898), .ZN(n708) );
  NAND2_X1 U761 ( .A1(n709), .A2(n708), .ZN(n717) );
  XNOR2_X1 U762 ( .A(G101), .B(n710), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n711), .B(KEYINPUT123), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U765 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U766 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U767 ( .A(KEYINPUT122), .B(n718), .ZN(G69) );
  XOR2_X1 U768 ( .A(n719), .B(KEYINPUT124), .Z(n720) );
  XNOR2_X1 U769 ( .A(n721), .B(n720), .ZN(n723) );
  XOR2_X1 U770 ( .A(n723), .B(n722), .Z(n727) );
  XNOR2_X1 U771 ( .A(n724), .B(n727), .ZN(n725) );
  NOR2_X1 U772 ( .A1(n725), .A2(G953), .ZN(n726) );
  XNOR2_X1 U773 ( .A(KEYINPUT125), .B(n726), .ZN(n731) );
  XNOR2_X1 U774 ( .A(n727), .B(G227), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U778 ( .A(G131), .B(KEYINPUT127), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(n732), .ZN(G33) );
  XNOR2_X1 U780 ( .A(G140), .B(n734), .ZN(G42) );
endmodule

