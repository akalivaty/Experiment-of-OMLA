

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n975), .ZN(n760) );
  INV_X1 U552 ( .A(n725), .ZN(n726) );
  AND2_X1 U553 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U554 ( .A1(n779), .A2(n760), .ZN(n761) );
  AND2_X1 U555 ( .A1(n578), .A2(n577), .ZN(n517) );
  XOR2_X1 U556 ( .A(KEYINPUT76), .B(n607), .Z(n518) );
  NOR2_X1 U557 ( .A1(n752), .A2(n749), .ZN(n730) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n716) );
  XNOR2_X1 U559 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n737) );
  NAND2_X1 U560 ( .A1(n726), .A2(G8), .ZN(n727) );
  XNOR2_X1 U561 ( .A(n727), .B(KEYINPUT91), .ZN(n768) );
  INV_X1 U562 ( .A(KEYINPUT17), .ZN(n560) );
  XNOR2_X1 U563 ( .A(n611), .B(KEYINPUT15), .ZN(n967) );
  NOR2_X1 U564 ( .A1(G543), .A2(n526), .ZN(n519) );
  XNOR2_X1 U565 ( .A(n561), .B(n560), .ZN(n888) );
  XOR2_X1 U566 ( .A(KEYINPUT67), .B(n521), .Z(n663) );
  XNOR2_X1 U567 ( .A(KEYINPUT75), .B(n603), .ZN(n971) );
  AND2_X1 U568 ( .A1(n888), .A2(G138), .ZN(n581) );
  INV_X1 U569 ( .A(G651), .ZN(n526) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n519), .Z(n654) );
  NAND2_X1 U571 ( .A1(G63), .A2(n654), .ZN(n523) );
  XNOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .ZN(n520) );
  XNOR2_X1 U573 ( .A(n520), .B(KEYINPUT69), .ZN(n642) );
  NOR2_X1 U574 ( .A1(n642), .A2(G651), .ZN(n521) );
  NAND2_X1 U575 ( .A1(G51), .A2(n663), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U577 ( .A(KEYINPUT6), .B(n524), .ZN(n532) );
  NOR2_X1 U578 ( .A1(G543), .A2(G651), .ZN(n655) );
  NAND2_X1 U579 ( .A1(n655), .A2(G89), .ZN(n525) );
  XNOR2_X1 U580 ( .A(n525), .B(KEYINPUT4), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n642), .A2(n526), .ZN(n658) );
  NAND2_X1 U582 ( .A1(G76), .A2(n658), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U584 ( .A(KEYINPUT77), .B(n529), .ZN(n530) );
  XNOR2_X1 U585 ( .A(KEYINPUT5), .B(n530), .ZN(n531) );
  NOR2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n534) );
  XOR2_X1 U587 ( .A(KEYINPUT78), .B(KEYINPUT7), .Z(n533) );
  XNOR2_X1 U588 ( .A(n534), .B(n533), .ZN(G168) );
  XNOR2_X1 U589 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n535) );
  XNOR2_X1 U590 ( .A(n535), .B(G168), .ZN(G286) );
  NAND2_X1 U591 ( .A1(G85), .A2(n655), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G72), .A2(n658), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G60), .A2(n654), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G47), .A2(n663), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U597 ( .A1(n541), .A2(n540), .ZN(G290) );
  XOR2_X1 U598 ( .A(G2443), .B(G2446), .Z(n543) );
  XNOR2_X1 U599 ( .A(G2427), .B(G2451), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n543), .B(n542), .ZN(n549) );
  XOR2_X1 U601 ( .A(G2430), .B(G2454), .Z(n545) );
  XNOR2_X1 U602 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U603 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U604 ( .A(G2435), .B(G2438), .Z(n546) );
  XNOR2_X1 U605 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U606 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U607 ( .A1(G14), .A2(n550), .ZN(G401) );
  XNOR2_X1 U608 ( .A(KEYINPUT71), .B(KEYINPUT9), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G90), .A2(n655), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G77), .A2(n658), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n554), .B(n553), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n654), .A2(G64), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n555), .B(KEYINPUT70), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G52), .A2(n663), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U619 ( .A1(G2104), .A2(G2105), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G135), .A2(n888), .ZN(n563) );
  AND2_X1 U621 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U622 ( .A1(G111), .A2(n892), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n570) );
  INV_X1 U624 ( .A(G2104), .ZN(n564) );
  NAND2_X1 U625 ( .A1(KEYINPUT68), .A2(n564), .ZN(n567) );
  INV_X1 U626 ( .A(KEYINPUT68), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n565), .A2(G2104), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n576) );
  INV_X1 U629 ( .A(G2105), .ZN(n574) );
  AND2_X1 U630 ( .A1(n576), .A2(G2105), .ZN(n586) );
  NAND2_X1 U631 ( .A1(n586), .A2(G123), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT18), .B(n568), .Z(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n572) );
  NOR2_X1 U634 ( .A1(n576), .A2(G2105), .ZN(n582) );
  BUF_X1 U635 ( .A(n582), .Z(n889) );
  NAND2_X1 U636 ( .A1(n889), .A2(G99), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n917) );
  XNOR2_X1 U638 ( .A(G2096), .B(n917), .ZN(n573) );
  OR2_X1 U639 ( .A1(G2100), .A2(n573), .ZN(G156) );
  NAND2_X1 U640 ( .A1(G126), .A2(n586), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G114), .A2(n892), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n574), .A2(G102), .ZN(n575) );
  OR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n579), .A2(n517), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(G164) );
  INV_X1 U646 ( .A(G57), .ZN(G237) );
  INV_X1 U647 ( .A(G132), .ZN(G219) );
  INV_X1 U648 ( .A(G82), .ZN(G220) );
  NAND2_X1 U649 ( .A1(n892), .A2(G113), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G101), .A2(n582), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT23), .B(n583), .Z(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G137), .A2(n888), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G125), .A2(n586), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U656 ( .A1(n590), .A2(n589), .ZN(G160) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n834) );
  NAND2_X1 U660 ( .A1(n834), .A2(G567), .ZN(n592) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n592), .Z(G234) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n594) );
  NAND2_X1 U663 ( .A1(G56), .A2(n654), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n594), .B(n593), .ZN(n602) );
  NAND2_X1 U665 ( .A1(n655), .A2(G81), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT12), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G68), .A2(n658), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT13), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G43), .A2(n663), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  INV_X1 U673 ( .A(n971), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n604), .A2(G860), .ZN(G153) );
  INV_X1 U675 ( .A(G171), .ZN(G301) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U677 ( .A1(G54), .A2(n663), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G92), .A2(n655), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G79), .A2(n658), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n654), .A2(G66), .ZN(n607) );
  NOR2_X1 U682 ( .A1(n608), .A2(n518), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U684 ( .A(n967), .ZN(n624) );
  INV_X1 U685 ( .A(G868), .ZN(n676) );
  NAND2_X1 U686 ( .A1(n624), .A2(n676), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U688 ( .A1(G78), .A2(n658), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G53), .A2(n663), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G65), .A2(n654), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G91), .A2(n655), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n620), .B(KEYINPUT72), .ZN(n977) );
  XNOR2_X1 U696 ( .A(KEYINPUT73), .B(n977), .ZN(G299) );
  NAND2_X1 U697 ( .A1(G868), .A2(G286), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G299), .A2(n676), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G297) );
  INV_X1 U700 ( .A(G559), .ZN(n626) );
  NOR2_X1 U701 ( .A1(G860), .A2(n626), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U703 ( .A(KEYINPUT16), .B(n625), .Z(G148) );
  NAND2_X1 U704 ( .A1(n626), .A2(n967), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n627), .A2(G868), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n971), .A2(n676), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G559), .A2(n967), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT80), .ZN(n673) );
  XOR2_X1 U710 ( .A(n673), .B(KEYINPUT81), .Z(n631) );
  XNOR2_X1 U711 ( .A(n971), .B(n631), .ZN(n632) );
  NOR2_X1 U712 ( .A1(G860), .A2(n632), .ZN(n633) );
  XOR2_X1 U713 ( .A(n633), .B(KEYINPUT82), .Z(n641) );
  NAND2_X1 U714 ( .A1(G67), .A2(n654), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G80), .A2(n658), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G93), .A2(n655), .ZN(n636) );
  XNOR2_X1 U718 ( .A(KEYINPUT83), .B(n636), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n663), .A2(G55), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n675) );
  XNOR2_X1 U722 ( .A(n641), .B(n675), .ZN(G145) );
  NAND2_X1 U723 ( .A1(G49), .A2(n663), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G87), .A2(n642), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U726 ( .A1(n654), .A2(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G651), .A2(G74), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G88), .A2(n655), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G75), .A2(n658), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G62), .A2(n654), .ZN(n651) );
  NAND2_X1 U733 ( .A1(G50), .A2(n663), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U735 ( .A1(n653), .A2(n652), .ZN(G166) );
  NAND2_X1 U736 ( .A1(G61), .A2(n654), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G86), .A2(n655), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n658), .A2(G73), .ZN(n659) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n659), .Z(n660) );
  NOR2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n662), .B(KEYINPUT84), .ZN(n665) );
  NAND2_X1 U743 ( .A1(G48), .A2(n663), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n665), .A2(n664), .ZN(G305) );
  XOR2_X1 U745 ( .A(G290), .B(G288), .Z(n666) );
  XNOR2_X1 U746 ( .A(n971), .B(n666), .ZN(n669) );
  XOR2_X1 U747 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n667) );
  XNOR2_X1 U748 ( .A(n675), .B(n667), .ZN(n668) );
  XOR2_X1 U749 ( .A(n669), .B(n668), .Z(n671) );
  XNOR2_X1 U750 ( .A(G166), .B(G299), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(G305), .ZN(n908) );
  XNOR2_X1 U753 ( .A(n673), .B(n908), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n674), .A2(G868), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U765 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U766 ( .A1(G96), .A2(n685), .ZN(n838) );
  NAND2_X1 U767 ( .A1(G2106), .A2(n838), .ZN(n689) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n686) );
  NOR2_X1 U769 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G108), .A2(n687), .ZN(n839) );
  NAND2_X1 U771 ( .A1(G567), .A2(n839), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n840) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n840), .A2(n690), .ZN(n837) );
  NAND2_X1 U775 ( .A1(n837), .A2(G36), .ZN(G176) );
  XOR2_X1 U776 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NOR2_X2 U777 ( .A1(G164), .A2(G1384), .ZN(n800) );
  XNOR2_X1 U778 ( .A(n800), .B(KEYINPUT65), .ZN(n692) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n801) );
  NOR2_X1 U780 ( .A1(n692), .A2(n801), .ZN(n725) );
  BUF_X1 U781 ( .A(n725), .Z(n718) );
  INV_X1 U782 ( .A(KEYINPUT93), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n718), .B(n693), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n695), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n694), .B(KEYINPUT27), .ZN(n697) );
  INV_X1 U786 ( .A(G1956), .ZN(n1002) );
  BUF_X1 U787 ( .A(n695), .Z(n720) );
  NOR2_X1 U788 ( .A1(n1002), .A2(n720), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n711) );
  NOR2_X1 U790 ( .A1(n711), .A2(n977), .ZN(n698) );
  XOR2_X1 U791 ( .A(n698), .B(KEYINPUT28), .Z(n715) );
  AND2_X1 U792 ( .A1(n718), .A2(G1996), .ZN(n700) );
  XOR2_X1 U793 ( .A(KEYINPUT66), .B(KEYINPUT26), .Z(n699) );
  XNOR2_X1 U794 ( .A(n700), .B(n699), .ZN(n702) );
  INV_X1 U795 ( .A(n718), .ZN(n729) );
  NAND2_X1 U796 ( .A1(n729), .A2(G1341), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n971), .A2(n703), .ZN(n708) );
  NAND2_X1 U799 ( .A1(n967), .A2(n708), .ZN(n707) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n720), .ZN(n705) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n729), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n710) );
  OR2_X1 U804 ( .A1(n967), .A2(n708), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n711), .A2(n977), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U809 ( .A(n717), .B(n716), .ZN(n724) );
  NOR2_X1 U810 ( .A1(n718), .A2(G1961), .ZN(n719) );
  XOR2_X1 U811 ( .A(KEYINPUT92), .B(n719), .Z(n722) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n953) );
  NAND2_X1 U813 ( .A1(n720), .A2(n953), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n734) );
  NAND2_X1 U815 ( .A1(n734), .A2(G171), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n740) );
  INV_X1 U817 ( .A(G1966), .ZN(n728) );
  AND2_X1 U818 ( .A1(n768), .A2(n728), .ZN(n752) );
  NOR2_X1 U819 ( .A1(n729), .A2(G2084), .ZN(n749) );
  NAND2_X1 U820 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U821 ( .A(n731), .B(KEYINPUT94), .ZN(n732) );
  XNOR2_X1 U822 ( .A(KEYINPUT30), .B(n732), .ZN(n733) );
  NOR2_X1 U823 ( .A1(G168), .A2(n733), .ZN(n736) );
  NOR2_X1 U824 ( .A1(G171), .A2(n734), .ZN(n735) );
  NOR2_X1 U825 ( .A1(n736), .A2(n735), .ZN(n738) );
  XNOR2_X1 U826 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n750) );
  NAND2_X1 U828 ( .A1(n750), .A2(G286), .ZN(n745) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n729), .ZN(n742) );
  INV_X1 U830 ( .A(n768), .ZN(n779) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n779), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(G303), .A2(n743), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U835 ( .A(n746), .B(KEYINPUT96), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n747), .A2(G8), .ZN(n748) );
  XNOR2_X1 U837 ( .A(n748), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U838 ( .A1(G8), .A2(n749), .ZN(n754) );
  INV_X1 U839 ( .A(n750), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n777) );
  NOR2_X1 U843 ( .A1(G303), .A2(G1971), .ZN(n758) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n757) );
  XOR2_X1 U845 ( .A(KEYINPUT97), .B(n757), .Z(n983) );
  NOR2_X1 U846 ( .A1(n758), .A2(n983), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n777), .A2(n759), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n975) );
  XNOR2_X1 U849 ( .A(n763), .B(KEYINPUT64), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XNOR2_X1 U851 ( .A(n764), .B(KEYINPUT24), .ZN(n765) );
  AND2_X1 U852 ( .A1(n765), .A2(n768), .ZN(n772) );
  OR2_X1 U853 ( .A1(KEYINPUT33), .A2(n772), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n774) );
  XNOR2_X1 U855 ( .A(G1981), .B(G305), .ZN(n987) );
  AND2_X1 U856 ( .A1(n983), .A2(KEYINPUT33), .ZN(n769) );
  AND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U858 ( .A1(n987), .A2(n770), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n782) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G8), .A2(n775), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U865 ( .A(KEYINPUT98), .B(n780), .Z(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n816) );
  NAND2_X1 U867 ( .A1(n586), .A2(G129), .ZN(n789) );
  NAND2_X1 U868 ( .A1(G141), .A2(n888), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G117), .A2(n892), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n889), .A2(G105), .ZN(n785) );
  XOR2_X1 U872 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U875 ( .A(KEYINPUT89), .B(n790), .Z(n902) );
  NAND2_X1 U876 ( .A1(G1996), .A2(n902), .ZN(n799) );
  NAND2_X1 U877 ( .A1(G131), .A2(n888), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G107), .A2(n892), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n586), .A2(G119), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT88), .B(n793), .Z(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n889), .A2(G95), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n878) );
  NAND2_X1 U885 ( .A1(G1991), .A2(n878), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n923) );
  XOR2_X1 U887 ( .A(n800), .B(KEYINPUT65), .Z(n802) );
  NOR2_X1 U888 ( .A1(n802), .A2(n801), .ZN(n829) );
  NAND2_X1 U889 ( .A1(n923), .A2(n829), .ZN(n803) );
  XOR2_X1 U890 ( .A(KEYINPUT90), .B(n803), .Z(n821) );
  INV_X1 U891 ( .A(n821), .ZN(n814) );
  XOR2_X1 U892 ( .A(KEYINPUT37), .B(G2067), .Z(n826) );
  NAND2_X1 U893 ( .A1(n888), .A2(G140), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT87), .B(n804), .Z(n806) );
  NAND2_X1 U895 ( .A1(n889), .A2(G104), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n807), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G128), .A2(n586), .ZN(n809) );
  NAND2_X1 U899 ( .A1(G116), .A2(n892), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  NOR2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U903 ( .A(KEYINPUT36), .B(n813), .Z(n899) );
  AND2_X1 U904 ( .A1(n826), .A2(n899), .ZN(n930) );
  NAND2_X1 U905 ( .A1(n829), .A2(n930), .ZN(n824) );
  NAND2_X1 U906 ( .A1(n814), .A2(n824), .ZN(n815) );
  NOR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n974) );
  NAND2_X1 U909 ( .A1(n974), .A2(n829), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n832) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n902), .ZN(n934) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n878), .ZN(n920) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n920), .A2(n819), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U916 ( .A1(n934), .A2(n822), .ZN(n823) );
  XNOR2_X1 U917 ( .A(KEYINPUT39), .B(n823), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n828) );
  NOR2_X1 U919 ( .A1(n826), .A2(n899), .ZN(n827) );
  XNOR2_X1 U920 ( .A(KEYINPUT99), .B(n827), .ZN(n939) );
  NAND2_X1 U921 ( .A1(n828), .A2(n939), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U924 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT100), .B(n840), .Z(G319) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n841), .B(KEYINPUT42), .ZN(n851) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(KEYINPUT102), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT101), .B(G2096), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(G2100), .B(G2084), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT103), .B(G2678), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U949 ( .A(KEYINPUT105), .B(G1956), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1961), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n854), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G1966), .B(G1971), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1981), .B(G1976), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT104), .B(G2474), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n889), .A2(G100), .ZN(n869) );
  NAND2_X1 U962 ( .A1(G136), .A2(n888), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G112), .A2(n892), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n586), .A2(G124), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT44), .B(n865), .Z(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT106), .B(n870), .Z(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT107), .B(KEYINPUT110), .Z(n872) );
  XNOR2_X1 U971 ( .A(G164), .B(KEYINPUT109), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT46), .B(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n917), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U976 ( .A(G160), .B(n876), .Z(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G130), .A2(n586), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G118), .A2(n892), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G142), .A2(n888), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G106), .A2(n889), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(n887), .B(n886), .Z(n901) );
  NAND2_X1 U987 ( .A1(G139), .A2(n888), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U990 ( .A1(n892), .A2(G115), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(KEYINPUT108), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G127), .A2(n586), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n924) );
  XNOR2_X1 U996 ( .A(n899), .B(n924), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U998 ( .A(n903), .B(n902), .Z(n904) );
  XNOR2_X1 U999 ( .A(G162), .B(n904), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(G286), .B(KEYINPUT111), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(G171), .B(n967), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n910), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n913), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n914), .B(KEYINPUT112), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n963) );
  XOR2_X1 U1016 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n942) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(KEYINPUT113), .B(n921), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n932) );
  XOR2_X1 U1022 ( .A(n924), .B(KEYINPUT115), .Z(n925) );
  XOR2_X1 U1023 ( .A(G2072), .B(n925), .Z(n927) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT50), .B(n928), .Z(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(KEYINPUT51), .B(n935), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT114), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n963), .A2(n943), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n944), .A2(G29), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(n945), .B(KEYINPUT118), .ZN(n998) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n958) );
  XNOR2_X1 U1040 ( .A(G1996), .B(G32), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n952) );
  XOR2_X1 U1043 ( .A(G2067), .B(G26), .Z(n948) );
  NAND2_X1 U1044 ( .A1(n948), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G25), .B(G1991), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1048 ( .A(G27), .B(n953), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1056 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n966), .A2(G11), .ZN(n996) );
  XOR2_X1 U1059 ( .A(KEYINPUT56), .B(G16), .Z(n994) );
  XNOR2_X1 U1060 ( .A(n967), .B(G1348), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G171), .B(G1961), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT119), .B(n970), .ZN(n982) );
  XNOR2_X1 U1064 ( .A(G1341), .B(KEYINPUT122), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n980) );
  XOR2_X1 U1068 ( .A(G1956), .B(n977), .Z(n978) );
  XNOR2_X1 U1069 ( .A(KEYINPUT120), .B(n978), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n992) );
  XOR2_X1 U1072 ( .A(n983), .B(KEYINPUT121), .Z(n985) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G303), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n990) );
  XOR2_X1 U1075 ( .A(G1966), .B(G168), .Z(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1077 ( .A(KEYINPUT57), .B(n988), .Z(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1082 ( .A1(n998), .A2(n997), .ZN(n1027) );
  XOR2_X1 U1083 ( .A(G1966), .B(G21), .Z(n1013) );
  XOR2_X1 U1084 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n999) );
  XNOR2_X1 U1085 ( .A(KEYINPUT60), .B(n999), .ZN(n1011) );
  XOR2_X1 U1086 ( .A(G4), .B(KEYINPUT124), .Z(n1001) );
  XNOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1001), .B(n1000), .ZN(n1009) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(n1002), .B(G20), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(KEYINPUT123), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1011), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(KEYINPUT127), .B(n1014), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(G1961), .B(G5), .Z(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1101 ( .A(G1976), .B(G23), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1025), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(n1028), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

