//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT13), .ZN(new_n203));
  INV_X1    g002(.A(G8gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G1gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n204), .B1(new_n206), .B2(KEYINPUT86), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(new_n208), .B2(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n207), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT14), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT15), .B(new_n212), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n215), .B(KEYINPUT85), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n212), .B(KEYINPUT15), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n211), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n211), .A2(new_n221), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n203), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n207), .B(new_n210), .Z(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n226), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(new_n202), .A3(new_n223), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n224), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n223), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT87), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT11), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT12), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n232), .B(new_n243), .C1(new_n235), .C2(new_n236), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT27), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G183gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253));
  AOI21_X1  g052(.A(G190gat), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT27), .B(G183gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n254), .B(new_n259), .C1(new_n253), .C2(new_n255), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(KEYINPUT28), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n268), .A2(new_n269), .B1(new_n267), .B2(new_n266), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT68), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n264), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n266), .B(KEYINPUT23), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G183gat), .B(G190gat), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .A4(new_n265), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n282), .A2(new_n283), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n265), .B2(KEYINPUT65), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(KEYINPUT65), .B2(new_n265), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n278), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n250), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT74), .B(G218gat), .Z(new_n296));
  OAI211_X1 g095(.A(G211gat), .B(new_n295), .C1(new_n296), .C2(KEYINPUT22), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G218gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n249), .B1(new_n278), .B2(new_n291), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n294), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n301), .B(G218gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n261), .A2(new_n263), .B1(new_n274), .B2(KEYINPUT69), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n290), .B1(new_n307), .B2(new_n277), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n249), .B1(new_n308), .B2(KEYINPUT29), .ZN(new_n309));
  INV_X1    g108(.A(new_n304), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT37), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT38), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n303), .B1(new_n294), .B2(new_n304), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n306), .A3(new_n310), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT37), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G8gat), .B(G36gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G64gat), .ZN(new_n319));
  INV_X1    g118(.A(G92gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n312), .A2(new_n313), .A3(new_n317), .A4(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n329), .B2(KEYINPUT2), .ZN(new_n330));
  XOR2_X1   g129(.A(G141gat), .B(G148gat), .Z(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(KEYINPUT2), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(new_n327), .A3(new_n328), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n336), .A2(new_n337), .B1(G155gat), .B2(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n337), .ZN(new_n341));
  NOR3_X1   g140(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n326), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(KEYINPUT76), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n332), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  INV_X1    g145(.A(G120gat), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT1), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n348), .B(new_n349), .C1(new_n346), .C2(new_n347), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n346), .A2(new_n347), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(G113gat), .B2(G120gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT70), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G127gat), .B(G134gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n351), .A2(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n349), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n332), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n343), .A2(KEYINPUT76), .B1(new_n331), .B2(new_n333), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n339), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n360), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n325), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT71), .A3(new_n359), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n366), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n376));
  NOR2_X1   g175(.A1(new_n345), .A2(new_n361), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n332), .C1(new_n340), .C2(new_n344), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n361), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n369), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n371), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(new_n325), .A3(new_n369), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G57gat), .ZN(new_n391));
  INV_X1    g190(.A(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n385), .A2(new_n387), .A3(new_n393), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n396), .B(new_n393), .C1(new_n385), .C2(new_n387), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n314), .A2(new_n315), .A3(new_n321), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT84), .B1(new_n324), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(new_n396), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n393), .B1(new_n385), .B2(new_n387), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n399), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n323), .A4(new_n401), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n312), .A2(new_n317), .A3(new_n322), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT38), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n369), .B1(new_n386), .B2(new_n383), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n362), .A2(new_n367), .A3(new_n369), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT39), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT82), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n419), .A3(KEYINPUT39), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n415), .B(new_n393), .C1(new_n421), .C2(new_n413), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n395), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT30), .A4(new_n321), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n322), .B1(new_n305), .B2(new_n311), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n321), .B1(new_n314), .B2(new_n315), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n430), .B2(new_n401), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n429), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G50gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G22gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(G228gat), .A2(G233gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n306), .A2(new_n293), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n366), .B1(new_n447), .B2(new_n381), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n382), .A2(new_n293), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n303), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n381), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n345), .ZN(new_n454));
  INV_X1    g253(.A(new_n446), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n450), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n445), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n444), .B1(new_n457), .B2(KEYINPUT80), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n448), .A2(new_n446), .A3(new_n451), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n455), .B1(new_n454), .B2(new_n450), .ZN(new_n460));
  OAI21_X1  g259(.A(G22gat), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n452), .A2(new_n445), .A3(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n461), .A2(KEYINPUT80), .A3(new_n462), .A4(new_n444), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n412), .A2(new_n440), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n373), .A2(new_n374), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n292), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n278), .A2(new_n374), .A3(new_n373), .A4(new_n291), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  NAND2_X1  g271(.A1(G227gat), .A2(G233gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT64), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n472), .B1(new_n471), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT72), .B(G71gat), .ZN(new_n479));
  INV_X1    g278(.A(G99gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G15gat), .B(G43gat), .Z(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n474), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n469), .B2(new_n470), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n485), .B2(KEYINPUT33), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT32), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI221_X4 g288(.A(new_n487), .B1(KEYINPUT33), .B2(new_n483), .C1(new_n471), .C2(new_n474), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n478), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n474), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(new_n483), .ZN(new_n496));
  INV_X1    g295(.A(new_n490), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n469), .A2(new_n470), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT34), .B1(new_n498), .B2(new_n484), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n475), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT36), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT73), .B1(new_n489), .B2(new_n490), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n491), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n478), .B(KEYINPUT73), .C1(new_n489), .C2(new_n490), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n502), .B1(new_n506), .B2(KEYINPUT36), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT78), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n407), .B2(new_n434), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n398), .A2(new_n400), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(new_n438), .A3(KEYINPUT78), .A4(new_n432), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n464), .A2(new_n465), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n467), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n504), .A2(new_n466), .A3(new_n505), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n513), .A2(KEYINPUT35), .A3(new_n407), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n435), .A2(new_n439), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n491), .A2(new_n501), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n248), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT21), .ZN(new_n524));
  NAND2_X1  g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT88), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  INV_X1    g329(.A(G57gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G64gat), .ZN(new_n532));
  INV_X1    g331(.A(G64gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G57gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n533), .B2(G57gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n531), .A2(KEYINPUT89), .A3(G64gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n534), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(new_n537), .A3(new_n530), .A4(new_n528), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n225), .B1(new_n524), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT92), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n551), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n549), .A2(new_n524), .ZN(new_n557));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT93), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(KEYINPUT7), .ZN(new_n571));
  AND2_X1   g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(KEYINPUT95), .A2(G99gat), .A3(G106gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n392), .A2(KEYINPUT96), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G85gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n585), .A3(new_n320), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n568), .B1(new_n576), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n572), .ZN(new_n589));
  INV_X1    g388(.A(new_n570), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n574), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT96), .B(G85gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n320), .A2(new_n594), .B1(new_n580), .B2(new_n581), .ZN(new_n595));
  INV_X1    g394(.A(new_n568), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(KEYINPUT97), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n599), .B(new_n568), .C1(new_n576), .C2(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n221), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n227), .A2(new_n228), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n567), .B(new_n602), .C1(new_n603), .C2(new_n601), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(KEYINPUT98), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(KEYINPUT98), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n566), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n604), .A2(KEYINPUT98), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(KEYINPUT98), .ZN(new_n609));
  INV_X1    g408(.A(new_n566), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n607), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n607), .B2(new_n611), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n564), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n588), .A2(new_n539), .A3(new_n597), .A4(new_n544), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n544), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT90), .B1(new_n539), .B2(new_n544), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT99), .B1(new_n601), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n549), .A2(new_n626), .A3(new_n600), .A4(new_n598), .ZN(new_n627));
  AOI211_X1 g426(.A(KEYINPUT10), .B(new_n621), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n549), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n601), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n619), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n621), .B1(new_n625), .B2(new_n627), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n634), .A2(KEYINPUT100), .A3(new_n619), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT100), .B1(new_n634), .B2(new_n619), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT101), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n633), .A2(new_n635), .A3(new_n643), .A4(new_n636), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n618), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n523), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n510), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n519), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  AND2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n652), .A2(KEYINPUT42), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(KEYINPUT42), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n653), .B(new_n654), .C1(new_n204), .C2(new_n650), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n647), .B2(new_n507), .ZN(new_n656));
  INV_X1    g455(.A(new_n520), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n647), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n647), .A2(new_n466), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NOR3_X1   g461(.A1(new_n564), .A2(new_n617), .A3(new_n645), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n523), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n664), .A2(G29gat), .A3(new_n510), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT45), .Z(new_n666));
  NOR3_X1   g465(.A1(new_n564), .A2(new_n248), .A3(new_n645), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n515), .A2(new_n522), .ZN(new_n669));
  INV_X1    g468(.A(new_n617), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI211_X1 g470(.A(KEYINPUT44), .B(new_n617), .C1(new_n515), .C2(new_n522), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G29gat), .B1(new_n673), .B2(new_n510), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n666), .A2(new_n674), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n664), .A2(G36gat), .A3(new_n519), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT46), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n673), .B2(new_n519), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  OAI21_X1  g478(.A(G43gat), .B1(new_n673), .B2(new_n507), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n664), .A2(G43gat), .A3(new_n657), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n682), .B2(new_n684), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(G1330gat));
  OAI21_X1  g487(.A(G50gat), .B1(new_n673), .B2(new_n466), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n466), .A2(G50gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n664), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g491(.A(new_n645), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n618), .A2(new_n247), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n669), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n510), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n531), .ZN(G1332gat));
  XOR2_X1   g496(.A(new_n695), .B(KEYINPUT103), .Z(new_n698));
  AOI21_X1  g497(.A(new_n519), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n703));
  OAI22_X1  g502(.A1(new_n702), .A2(new_n703), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n703), .ZN(new_n705));
  NOR2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(G1333gat));
  NOR3_X1   g507(.A1(new_n695), .A2(G71gat), .A3(new_n657), .ZN(new_n709));
  INV_X1    g508(.A(new_n507), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n698), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(G71gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n513), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g514(.A1(new_n564), .A2(new_n693), .A3(new_n247), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n671), .B2(new_n672), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(KEYINPUT105), .B(new_n716), .C1(new_n671), .C2(new_n672), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n719), .A2(new_n407), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n617), .B1(new_n515), .B2(new_n522), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n564), .A2(new_n247), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(KEYINPUT51), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n645), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n407), .A2(new_n594), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n721), .A2(new_n594), .B1(new_n729), .B2(new_n730), .ZN(G1336gat));
  OAI21_X1  g530(.A(G92gat), .B1(new_n717), .B2(new_n519), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  INV_X1    g532(.A(new_n519), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n320), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n732), .B(new_n733), .C1(new_n729), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n734), .A3(new_n720), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n726), .A2(KEYINPUT106), .A3(new_n727), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n739), .A3(new_n725), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n735), .A2(new_n693), .ZN(new_n742));
  AOI22_X1  g541(.A1(G92gat), .A2(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n736), .B1(new_n743), .B2(new_n733), .ZN(G1337gat));
  OAI21_X1  g543(.A(new_n480), .B1(new_n729), .B2(new_n657), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n719), .A2(G99gat), .A3(new_n710), .A4(new_n720), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n719), .A2(new_n513), .A3(new_n720), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT107), .B(G106gat), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n466), .A2(new_n693), .A3(G106gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n740), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n738), .A2(new_n740), .A3(new_n751), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n750), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT53), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT53), .B1(new_n728), .B2(new_n751), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n749), .B1(new_n717), .B2(new_n466), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1339gat));
  NAND2_X1  g560(.A1(new_n646), .A2(new_n248), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n619), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n625), .A2(new_n627), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n629), .A3(new_n620), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(new_n766), .B2(new_n631), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n643), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n764), .A3(new_n631), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n771), .A3(KEYINPUT55), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n644), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n770), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n641), .B1(new_n633), .B2(KEYINPUT54), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT55), .B1(new_n769), .B2(new_n771), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n773), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n222), .A2(new_n223), .A3(new_n203), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n202), .B1(new_n229), .B2(new_n223), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n242), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n246), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n670), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n645), .A2(new_n786), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n782), .B2(new_n247), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n790), .B2(new_n670), .ZN(new_n791));
  INV_X1    g590(.A(new_n564), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n763), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n510), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n734), .A2(new_n516), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n247), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n772), .A2(new_n644), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n778), .B(KEYINPUT55), .C1(new_n769), .C2(new_n771), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n799), .B(new_n247), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n670), .B1(new_n802), .B2(new_n788), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n786), .B1(new_n615), .B2(new_n616), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n773), .B(new_n804), .C1(new_n779), .C2(new_n781), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n792), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n762), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n657), .A2(new_n513), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(new_n510), .A3(new_n734), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n248), .A2(new_n346), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n798), .B1(new_n810), .B2(new_n811), .ZN(G1340gat));
  OAI21_X1  g611(.A(new_n347), .B1(new_n796), .B2(new_n693), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(G120gat), .A3(new_n645), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT110), .Z(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n797), .A2(new_n817), .A3(new_n564), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n810), .A2(new_n564), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n817), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n617), .A2(G134gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n794), .A2(new_n795), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT56), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n734), .A2(new_n510), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n670), .A3(new_n824), .A4(new_n808), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n825), .A2(new_n826), .A3(G134gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n825), .B2(G134gat), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n823), .A2(KEYINPUT112), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n823), .B2(new_n829), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1343gat));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n833), .B(new_n834), .C1(new_n793), .C2(new_n466), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n466), .B1(new_n806), .B2(new_n762), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT113), .B1(new_n836), .B2(KEYINPUT57), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n466), .A2(new_n834), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n248), .A2(new_n780), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n789), .B1(new_n799), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n787), .B1(new_n840), .B2(new_n670), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n792), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n763), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n835), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n507), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n247), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G141gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n710), .A2(new_n466), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n248), .A2(G141gat), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n519), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n794), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT114), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT58), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n807), .A2(new_n407), .A3(new_n849), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n807), .A2(KEYINPUT115), .A3(new_n407), .A4(new_n849), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n519), .A3(new_n850), .A4(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n848), .A2(new_n856), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n856), .B1(new_n848), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(G1344gat));
  AOI21_X1  g665(.A(new_n693), .B1(new_n846), .B2(KEYINPUT118), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(KEYINPUT118), .B2(new_n846), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n763), .B1(new_n841), .B2(new_n792), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n834), .B1(new_n869), .B2(new_n466), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n807), .A2(new_n838), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G148gat), .B1(new_n872), .B2(KEYINPUT119), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT59), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n844), .A2(new_n846), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n693), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n859), .A2(new_n519), .A3(new_n860), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n877), .A3(new_n645), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1345gat));
  OAI21_X1  g683(.A(G155gat), .B1(new_n879), .B2(new_n792), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n327), .A3(new_n564), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1346gat));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n328), .A3(new_n670), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n879), .A2(new_n617), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(KEYINPUT120), .ZN(new_n890));
  OAI21_X1  g689(.A(G162gat), .B1(new_n889), .B2(KEYINPUT120), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1347gat));
  INV_X1    g691(.A(new_n516), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n519), .A2(new_n407), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n807), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n247), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n809), .A2(new_n407), .A3(new_n519), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n248), .A2(new_n240), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1348gat));
  INV_X1    g699(.A(G176gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n901), .A3(new_n645), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n898), .A2(new_n645), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n901), .ZN(G1349gat));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n807), .A2(new_n564), .A3(new_n808), .A4(new_n894), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G183gat), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n564), .A2(new_n255), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n895), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n910), .B2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n907), .B(new_n913), .C1(new_n895), .C2(new_n909), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n912), .B1(new_n911), .B2(new_n914), .ZN(new_n916));
  XNOR2_X1  g715(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n915), .A2(new_n916), .B1(new_n910), .B2(new_n917), .ZN(G1350gat));
  AOI21_X1  g717(.A(new_n262), .B1(new_n898), .B2(new_n670), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT61), .Z(new_n920));
  NAND3_X1  g719(.A1(new_n896), .A2(new_n262), .A3(new_n670), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n507), .A2(new_n894), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT124), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(new_n870), .B2(new_n871), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(G197gat), .A3(new_n247), .ZN(new_n926));
  INV_X1    g725(.A(new_n923), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n836), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n928), .A2(new_n247), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(G197gat), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n932), .A3(new_n645), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT126), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n925), .B2(new_n645), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(KEYINPUT62), .B2(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n928), .A2(new_n299), .A3(new_n564), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n925), .A2(new_n564), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n928), .B2(new_n670), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n670), .A2(new_n296), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT127), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n925), .B2(new_n946), .ZN(G1355gat));
endmodule


