//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n589, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G112), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n473), .B1(new_n476), .B2(G136), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n461), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(G162));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n462), .B2(new_n463), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n485), .B(new_n488), .C1(new_n463), .C2(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n490), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n491), .B1(new_n490), .B2(new_n497), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n502), .A2(G62), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT72), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n503), .B2(KEYINPUT71), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n501), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(G543), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n502), .A3(new_n515), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n509), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n508), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT5), .B(G543), .Z(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n501), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n524), .A2(G63), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n522), .B(new_n528), .C1(new_n529), .C2(new_n517), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  INV_X1    g106(.A(new_n517), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n501), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n501), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT73), .ZN(new_n541));
  AOI22_X1  g116(.A1(G43), .A2(new_n521), .B1(new_n532), .B2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OR3_X1    g125(.A1(new_n516), .A2(KEYINPUT9), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT9), .B1(new_n516), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n501), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n532), .B2(G91), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G166), .ZN(G303));
  INV_X1    g133(.A(G49), .ZN(new_n559));
  INV_X1    g134(.A(G87), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n559), .A2(new_n516), .B1(new_n517), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(G288));
  NAND2_X1  g140(.A1(new_n521), .A2(G48), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n501), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n514), .A2(G86), .A3(new_n502), .A4(new_n515), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(G47), .A2(new_n521), .B1(new_n532), .B2(G85), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT75), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n501), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n532), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT10), .Z(new_n578));
  NAND2_X1  g153(.A1(G79), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G66), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n523), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n521), .A2(G54), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n576), .B1(new_n584), .B2(G868), .ZN(G284));
  OAI21_X1  g160(.A(new_n576), .B1(new_n584), .B2(G868), .ZN(G321));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G286), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(G299), .B(KEYINPUT76), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n587), .ZN(G297));
  AOI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n587), .ZN(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n543), .A2(new_n587), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n583), .A2(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n587), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g172(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT12), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT13), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT77), .B(G2100), .Z(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  INV_X1    g178(.A(G111), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n604), .A2(KEYINPUT80), .A3(G2105), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT80), .B1(new_n604), .B2(G2105), .ZN(new_n606));
  OAI21_X1  g181(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n605), .A2(new_n608), .B1(new_n476), .B2(G135), .ZN(new_n609));
  INV_X1    g184(.A(G123), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n479), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n600), .A2(new_n601), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT79), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n603), .A2(new_n612), .A3(new_n614), .ZN(G156));
  INV_X1    g190(.A(G14), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT15), .B(G2435), .Z(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(G2438), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2427), .B(G2430), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n619), .A2(new_n622), .A3(new_n620), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT82), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT83), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n632), .A2(new_n637), .A3(new_n634), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n616), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n630), .A2(new_n631), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n630), .A2(new_n631), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n633), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n639), .A2(new_n643), .ZN(G401));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  INV_X1    g250(.A(G29), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G25), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n478), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G119), .ZN(new_n680));
  OAI21_X1  g255(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n681));
  INV_X1    g256(.A(G107), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G2105), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n476), .B2(G131), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n677), .B1(new_n686), .B2(new_n676), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(G290), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(G290), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(G24), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1986), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(G1986), .A3(new_n694), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n689), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(G16), .B1(new_n508), .B2(new_n519), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n690), .A2(G22), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT88), .Z(new_n703));
  AND3_X1   g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n700), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(G288), .A2(KEYINPUT87), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n562), .A2(new_n708), .A3(new_n564), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n709), .A3(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G23), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n566), .A2(new_n568), .A3(G16), .A4(new_n569), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n717));
  OR2_X1    g292(.A1(G6), .A2(G16), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(new_n721));
  OAI21_X1  g296(.A(G1981), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G1981), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n723), .A2(new_n724), .A3(new_n719), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n710), .A2(new_n712), .ZN(new_n727));
  INV_X1    g302(.A(new_n711), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n714), .A2(new_n715), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n726), .A2(new_n729), .A3(new_n713), .A4(new_n706), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT86), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n730), .B2(new_n732), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n699), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT89), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n699), .B(new_n738), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n737), .A2(KEYINPUT36), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT36), .B1(new_n737), .B2(new_n739), .ZN(new_n742));
  NOR2_X1   g317(.A1(G164), .A2(new_n676), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G27), .B2(new_n676), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT99), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT98), .B(G2078), .Z(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(new_n747), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G33), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT25), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n476), .A2(G139), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT3), .B(G2104), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G127), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n461), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n751), .B1(new_n762), .B2(new_n676), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2072), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT24), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n676), .B1(new_n765), .B2(G34), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G160), .B2(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G2084), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT94), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n676), .A2(G32), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT26), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n773), .B(new_n775), .C1(G141), .C2(new_n476), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n679), .A2(G129), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n772), .B1(new_n778), .B2(new_n676), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n764), .B(new_n769), .C1(new_n771), .C2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n690), .A2(G5), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G301), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT97), .Z(new_n787));
  NAND4_X1  g362(.A1(new_n748), .A2(new_n749), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G29), .A2(G35), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G162), .B2(G29), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT29), .B(G2090), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n690), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT23), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT100), .B(G1956), .Z(new_n797));
  XOR2_X1   g372(.A(new_n796), .B(new_n797), .Z(new_n798));
  AND2_X1   g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n690), .A2(G19), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT91), .Z(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n543), .B2(G16), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT92), .B(G1341), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n676), .A2(G26), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT28), .Z(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(G116), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(G2105), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n476), .B2(G140), .ZN(new_n812));
  INV_X1    g387(.A(G128), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n479), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n690), .A2(G21), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G286), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G1966), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n818), .A2(new_n819), .B1(new_n784), .B2(new_n785), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n806), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n779), .A2(new_n771), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G2084), .B2(new_n768), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n803), .A2(new_n805), .B1(new_n819), .B2(new_n818), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT30), .B(G28), .ZN(new_n825));
  OR2_X1    g400(.A1(KEYINPUT31), .A2(G11), .ZN(new_n826));
  NAND2_X1  g401(.A1(KEYINPUT31), .A2(G11), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n825), .A2(new_n676), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n611), .B2(new_n676), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT96), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n821), .A2(new_n823), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n690), .B1(new_n578), .B2(new_n582), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n690), .A2(G4), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT90), .B(G1348), .Z(new_n834));
  OR3_X1    g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n835), .A2(new_n836), .B1(new_n780), .B2(new_n781), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n799), .A2(new_n831), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n789), .A2(KEYINPUT101), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT101), .B1(new_n789), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n741), .A2(new_n742), .A3(new_n842), .ZN(G311));
  INV_X1    g418(.A(new_n742), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n740), .ZN(G150));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n532), .A2(G93), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n521), .A2(G55), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n848), .B(new_n849), .C1(new_n501), .C2(new_n850), .ZN(new_n851));
  OR3_X1    g426(.A1(new_n543), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n851), .A2(new_n847), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n847), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n543), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n583), .A2(new_n592), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n858), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n851), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(G145));
  NAND2_X1  g447(.A1(new_n776), .A2(new_n777), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n814), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n492), .A2(new_n496), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n487), .B2(new_n489), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n874), .A2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n762), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n476), .A2(G142), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n461), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n679), .B2(G130), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n599), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n685), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n778), .B(new_n814), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n490), .A2(new_n497), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n761), .A3(new_n877), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n880), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n611), .B(G160), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G162), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n880), .A2(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(new_n887), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n892), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n880), .A2(new_n902), .A3(new_n887), .A4(new_n891), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n903), .A2(new_n894), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n901), .B2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g485(.A(new_n856), .B(new_n595), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n583), .A2(G299), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n578), .A2(new_n553), .A3(new_n556), .A4(new_n582), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n915), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n921));
  INV_X1    g496(.A(G290), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(G303), .ZN(new_n923));
  NOR2_X1   g498(.A1(G290), .A2(G166), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n707), .A2(new_n709), .A3(G305), .ZN(new_n925));
  AOI21_X1  g500(.A(G305), .B1(new_n707), .B2(new_n709), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(G303), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(KEYINPUT106), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n916), .A2(new_n933), .A3(new_n919), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n921), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n921), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n851), .A2(new_n587), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  XNOR2_X1  g516(.A(G171), .B(G286), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n852), .B2(new_n855), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n852), .A2(new_n855), .A3(new_n942), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(new_n913), .A3(new_n914), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n945), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n943), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n918), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n931), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n931), .B(new_n946), .C1(new_n918), .C2(new_n948), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT108), .B(new_n941), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n952), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(KEYINPUT43), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT107), .B1(new_n957), .B2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n951), .A2(new_n961), .A3(new_n941), .A4(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n941), .B1(new_n951), .B2(new_n952), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n959), .A2(new_n963), .B1(new_n966), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n876), .B2(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(G160), .A2(G40), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n873), .B(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n814), .B(G2067), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n686), .A2(new_n688), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n686), .A2(new_n688), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n922), .A2(new_n696), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n922), .A2(new_n696), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n971), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n466), .A2(new_n469), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n968), .A2(G1384), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n876), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n498), .B2(new_n499), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(new_n968), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT56), .B(G2072), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n489), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n488), .B1(new_n757), .B2(new_n485), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT69), .B1(new_n998), .B2(new_n875), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n490), .A2(new_n491), .A3(new_n497), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n970), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT110), .B1(new_n889), .B2(new_n990), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1005), .B(G1384), .C1(new_n490), .C2(new_n497), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT50), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1956), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n984), .B1(new_n995), .B2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1002), .B(new_n990), .C1(new_n498), .C2(new_n499), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n986), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1956), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1011), .A2(new_n1012), .B1(new_n992), .B2(new_n993), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT116), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n553), .B2(new_n556), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1009), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1005), .B1(new_n876), .B2(G1384), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT110), .B(new_n990), .C1(new_n998), .C2(new_n875), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1002), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(new_n986), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(KEYINPUT115), .A3(new_n986), .A4(new_n1024), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n834), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1022), .A2(new_n986), .A3(new_n1023), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(G2067), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n583), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT114), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1010), .A2(new_n986), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1002), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1012), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND4_X1   g612(.A1(KEYINPUT114), .A2(new_n1037), .A3(new_n1018), .A4(new_n994), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n1021), .A2(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT61), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT118), .B(new_n1019), .C1(new_n995), .C2(new_n1008), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n1032), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n584), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1037), .A2(new_n1018), .A3(new_n994), .A4(KEYINPUT119), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1053), .A2(KEYINPUT61), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1020), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n989), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n972), .C1(new_n1001), .C2(KEYINPUT45), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n1031), .A2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1060), .A2(KEYINPUT117), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n544), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT59), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n544), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n583), .A4(new_n1032), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1058), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1039), .B1(new_n1052), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n987), .B1(new_n498), .B2(new_n499), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n986), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n819), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n970), .A2(G2084), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1028), .A2(new_n1024), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  NAND3_X1  g656(.A1(G286), .A2(new_n1081), .A3(G8), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(G286), .B2(G8), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT51), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(KEYINPUT122), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT121), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G286), .A2(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT120), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1082), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1089), .B2(new_n1085), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1087), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1092), .A2(new_n1082), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1079), .A2(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1027), .A2(new_n785), .A3(new_n1029), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n1104));
  OR4_X1    g679(.A1(new_n1104), .A2(new_n1074), .A3(G2078), .A4(new_n1075), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1059), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT109), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n991), .A2(new_n968), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n1059), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(G171), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1109), .B2(new_n1059), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT109), .B(new_n989), .C1(new_n991), .C2(new_n968), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1104), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n969), .A4(new_n1113), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT123), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(G301), .A3(new_n1103), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT54), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1108), .A2(new_n701), .A3(new_n1111), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1025), .A2(G2090), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1088), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G166), .A2(new_n1088), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1031), .A2(G8), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n724), .B1(new_n568), .B2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1133), .A2(G305), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(G305), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT49), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1131), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(KEYINPUT49), .A3(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n707), .A2(new_n709), .A3(G1976), .ZN(new_n1141));
  INV_X1    g716(.A(G1976), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT52), .B1(G288), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1141), .A2(new_n1143), .A3(G8), .A4(new_n1031), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(G8), .A3(new_n1031), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT52), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1140), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1011), .A2(G2090), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1088), .B1(new_n1124), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1130), .B(new_n1147), .C1(new_n1149), .C2(new_n1129), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1102), .A2(new_n1123), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n1152));
  AOI21_X1  g727(.A(G2078), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1103), .B(new_n1105), .C1(new_n1153), .C2(KEYINPUT53), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(new_n1154), .B2(G171), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(KEYINPUT124), .A3(G301), .A4(new_n1119), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1103), .A2(new_n1121), .ZN(new_n1159));
  OAI21_X1  g734(.A(G171), .B1(new_n1159), .B2(new_n1114), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1158), .B(KEYINPUT54), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1072), .A2(new_n1151), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1089), .A2(G168), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1150), .B2(new_n1167), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1166), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1169), .A2(new_n1130), .A3(new_n1147), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1150), .A2(new_n1115), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1099), .A2(new_n1101), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT62), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G288), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1140), .A2(new_n1142), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(G1981), .B2(G305), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1181), .A2(KEYINPUT113), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1131), .B1(new_n1181), .B2(KEYINPUT113), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1130), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1182), .A2(new_n1183), .B1(new_n1184), .B2(new_n1147), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1172), .A2(new_n1178), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n983), .B1(new_n1165), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n971), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n979), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n980), .A2(new_n1188), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(KEYINPUT48), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(KEYINPUT48), .B2(new_n1190), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n977), .B1(new_n975), .B2(new_n971), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n814), .A2(G2067), .ZN(new_n1194));
  OR3_X1    g769(.A1(new_n1193), .A2(KEYINPUT126), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT126), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1195), .A2(new_n971), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1188), .B1(new_n974), .B2(new_n778), .ZN(new_n1198));
  OR3_X1    g773(.A1(new_n1188), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT46), .B1(new_n1188), .B2(G1996), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n1192), .A2(new_n1197), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1187), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g780(.A1(G227), .A2(new_n459), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n674), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n639), .B2(new_n643), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1209), .A2(new_n909), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1210), .A2(new_n966), .ZN(G308));
  OAI211_X1 g785(.A(new_n1209), .B(new_n909), .C1(new_n965), .C2(new_n964), .ZN(G225));
endmodule


