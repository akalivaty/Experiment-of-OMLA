//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1320, new_n1321, new_n1322;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G238), .A3(G236), .A4(G237), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n453), .A2(KEYINPUT67), .A3(G567), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G125), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(new_n468), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n468), .A2(new_n464), .A3(G137), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n477), .A2(new_n480), .A3(new_n481), .ZN(G160));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n464), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(KEYINPUT70), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT71), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n475), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n468), .B1(new_n484), .B2(new_n487), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G124), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n478), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n500), .B(new_n501), .C1(new_n470), .C2(new_n471), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT72), .A2(G114), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT72), .A2(G114), .ZN(new_n506));
  OAI21_X1  g081(.A(G2105), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(G126), .A2(G2105), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n509), .B1(new_n464), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n468), .A2(new_n464), .A3(KEYINPUT4), .A4(G138), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n504), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(new_n519), .B1(new_n516), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT75), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n521), .B1(new_n520), .B2(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(KEYINPUT76), .B(G651), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  OR2_X1    g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n518), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G50), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT6), .B(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G88), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n529), .A2(new_n530), .A3(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT77), .B1(new_n520), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n548));
  AOI22_X1  g123(.A1(G51), .A2(new_n533), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G89), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n536), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n545), .A2(new_n551), .ZN(G168));
  AOI22_X1  g127(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G651), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT78), .B(G52), .Z(new_n556));
  NAND2_X1  g131(.A1(new_n533), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n536), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n555), .A2(new_n559), .ZN(G171));
  NAND2_X1  g135(.A1(new_n520), .A2(G56), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n554), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n520), .A2(G81), .A3(new_n535), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n533), .A2(G43), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n517), .A2(new_n519), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n516), .A2(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(G65), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  AND2_X1   g153(.A1(KEYINPUT6), .A2(G651), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT6), .A2(G651), .ZN(new_n580));
  OAI211_X1 g155(.A(G53), .B(G543), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(KEYINPUT79), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n535), .A2(G53), .A3(new_n583), .A4(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n520), .A2(G91), .A3(new_n535), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n578), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(G299));
  OAI221_X1 g167(.A(new_n557), .B1(new_n536), .B2(new_n558), .C1(new_n553), .C2(new_n554), .ZN(G301));
  INV_X1    g168(.A(G168), .ZN(G286));
  NAND3_X1  g169(.A1(new_n520), .A2(G87), .A3(new_n535), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n533), .A2(G49), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(KEYINPUT81), .B(G651), .C1(new_n520), .C2(G74), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G288));
  NAND3_X1  g178(.A1(new_n573), .A2(G61), .A3(new_n574), .ZN(new_n604));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n520), .A2(G86), .A3(new_n535), .ZN(new_n608));
  OAI211_X1 g183(.A(G48), .B(G543), .C1(new_n579), .C2(new_n580), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n554), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n533), .A2(G47), .ZN(new_n615));
  INV_X1    g190(.A(G85), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n536), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n520), .A2(G66), .ZN(new_n621));
  INV_X1    g196(.A(G79), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n518), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n573), .A2(G92), .A3(new_n574), .A4(new_n535), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT83), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n520), .A2(new_n628), .A3(G92), .A4(new_n535), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n626), .B2(new_n629), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n620), .B1(new_n633), .B2(G868), .ZN(G284));
  OAI21_X1  g209(.A(new_n620), .B1(new_n633), .B2(G868), .ZN(G321));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(G299), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(G168), .ZN(G297));
  OAI21_X1  g213(.A(new_n637), .B1(new_n636), .B2(G168), .ZN(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n633), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n633), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n464), .A2(new_n479), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT13), .Z(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(KEYINPUT84), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(KEYINPUT84), .ZN(new_n651));
  MUX2_X1   g226(.A(new_n650), .B(new_n648), .S(new_n651), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n488), .A2(G135), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT85), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  INV_X1    g230(.A(G111), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n655), .B1(new_n475), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n494), .B2(G123), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(G2096), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(G2096), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n652), .A2(new_n660), .A3(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2438), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2427), .B(G2430), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT14), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n673), .B1(new_n668), .B2(new_n671), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n668), .A2(new_n671), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n665), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AOI211_X1 g255(.A(new_n678), .B(new_n664), .C1(new_n674), .C2(new_n676), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n663), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2451), .B(G2454), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT16), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(new_n664), .ZN(new_n688));
  INV_X1    g263(.A(new_n663), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n677), .A2(new_n679), .A3(new_n665), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n682), .A2(new_n684), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G14), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n684), .B1(new_n682), .B2(new_n691), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT88), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n682), .A2(new_n691), .ZN(new_n696));
  INV_X1    g271(.A(new_n684), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n698), .A2(new_n699), .A3(G14), .A4(new_n692), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G401));
  XNOR2_X1  g277(.A(G2067), .B(G2678), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G2072), .A2(G2078), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n442), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G2084), .B(G2090), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT18), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n707), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n707), .B(KEYINPUT17), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n711), .B(new_n708), .C1(new_n705), .C2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n708), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(new_n705), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(G2096), .B(G2100), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G227));
  XNOR2_X1  g293(.A(G1981), .B(G1986), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1971), .B(G1976), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT19), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(G1956), .B(G2474), .Z(new_n724));
  XOR2_X1   g299(.A(G1961), .B(G1966), .Z(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n724), .A2(new_n725), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(new_n731), .B(new_n730), .S(new_n723), .Z(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(G1991), .B(G1996), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n733), .B(new_n734), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n737), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n720), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n737), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n736), .A2(new_n738), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(new_n744), .A3(new_n719), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n742), .A2(new_n745), .ZN(G229));
  INV_X1    g321(.A(KEYINPUT98), .ZN(new_n747));
  NOR2_X1   g322(.A1(G6), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT82), .B1(new_n533), .B2(G48), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n609), .A2(new_n610), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n608), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n554), .B1(new_n604), .B2(new_n605), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n748), .B1(new_n753), .B2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT32), .B(G1981), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT90), .Z(new_n757));
  INV_X1    g332(.A(G16), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G23), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n602), .B2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT33), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1976), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G22), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G166), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G1971), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n757), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT34), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(KEYINPUT34), .ZN(new_n769));
  INV_X1    g344(.A(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G25), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n488), .A2(G131), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n494), .A2(G119), .ZN(new_n773));
  OAI221_X1 g348(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(new_n770), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT35), .B(G1991), .Z(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n777), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n758), .A2(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n618), .B2(new_n758), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n768), .A2(new_n769), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT36), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n768), .A2(new_n787), .A3(new_n769), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n770), .A2(G35), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT95), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n496), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n792), .B(KEYINPUT97), .ZN(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n795), .A2(new_n798), .A3(new_n800), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n758), .A2(G4), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n633), .B2(new_n758), .ZN(new_n806));
  INV_X1    g381(.A(G1348), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n488), .A2(G141), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n494), .A2(G129), .ZN(new_n810));
  NAND3_X1  g385(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT26), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n813), .A2(new_n814), .B1(G105), .B2(new_n479), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n770), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n770), .B2(G32), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT27), .B(G1996), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT93), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT24), .ZN(new_n822));
  INV_X1    g397(.A(G34), .ZN(new_n823));
  AOI21_X1  g398(.A(G29), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G160), .B2(new_n770), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n818), .A2(new_n819), .B1(G2084), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(G301), .A2(G16), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n758), .A2(G5), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(G1961), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n758), .A2(G20), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT23), .ZN(new_n834));
  INV_X1    g409(.A(G299), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n758), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1956), .Z(new_n837));
  NAND3_X1  g412(.A1(new_n821), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT25), .ZN(new_n839));
  NAND2_X1  g414(.A1(G103), .A2(G2104), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n475), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n464), .A2(G127), .ZN(new_n843));
  NAND2_X1  g418(.A1(G115), .A2(G2104), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n841), .A2(new_n842), .B1(new_n845), .B2(new_n475), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n488), .A2(G139), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G29), .ZN(new_n851));
  NOR2_X1   g426(.A1(G29), .A2(G33), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT91), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G2072), .ZN(new_n855));
  NAND2_X1  g430(.A1(G164), .A2(G29), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G27), .B2(G29), .ZN(new_n857));
  INV_X1    g432(.A(G2078), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n659), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G29), .ZN(new_n861));
  INV_X1    g436(.A(G28), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT30), .ZN(new_n863));
  AOI21_X1  g438(.A(G29), .B1(new_n862), .B2(KEYINPUT30), .ZN(new_n864));
  OR2_X1    g439(.A1(KEYINPUT31), .A2(G11), .ZN(new_n865));
  NAND2_X1  g440(.A1(KEYINPUT31), .A2(G11), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n863), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n857), .A2(new_n858), .ZN(new_n868));
  AND4_X1   g443(.A1(new_n859), .A2(new_n861), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G1961), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n830), .A2(new_n870), .B1(new_n826), .B2(G2084), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n758), .A2(G19), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n567), .B2(new_n758), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(G1341), .Z(new_n874));
  NAND4_X1  g449(.A1(new_n855), .A2(new_n869), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n758), .A2(G21), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G168), .B2(new_n758), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT94), .B(G1966), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n770), .A2(G26), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT28), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n484), .A2(new_n487), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(G140), .A3(new_n478), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(G128), .A3(new_n475), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n885));
  INV_X1    g460(.A(G116), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n475), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n881), .B1(new_n890), .B2(new_n770), .ZN(new_n891));
  INV_X1    g466(.A(G2067), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n879), .B(new_n893), .C1(new_n854), .C2(G2072), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n838), .A2(new_n875), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n804), .A2(new_n808), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n747), .B1(new_n789), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g473(.A(KEYINPUT98), .B(new_n896), .C1(new_n786), .C2(new_n788), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G311));
  NAND2_X1  g475(.A1(new_n789), .A2(new_n897), .ZN(G150));
  NAND2_X1  g476(.A1(new_n633), .A2(G559), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n561), .A2(new_n562), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G651), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n564), .A2(new_n565), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n520), .A2(G93), .A3(new_n535), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n533), .A2(G55), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n573), .A2(G67), .A3(new_n574), .ZN(new_n910));
  NAND2_X1  g485(.A1(G80), .A2(G543), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G651), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n905), .A2(new_n906), .A3(new_n909), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(new_n908), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n554), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n563), .A2(new_n566), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n903), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT39), .ZN(new_n920));
  AOI21_X1  g495(.A(G860), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(G860), .B1(new_n915), .B2(new_n916), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT37), .Z(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT99), .Z(G145));
  OR2_X1    g501(.A1(new_n496), .A2(G160), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n496), .A2(G160), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n860), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n860), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n935));
  INV_X1    g510(.A(G118), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n475), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n488), .B2(G142), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n494), .A2(KEYINPUT100), .A3(G130), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT100), .B1(new_n494), .B2(G130), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n647), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n647), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n943), .A2(new_n775), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n775), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n934), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n889), .A2(G164), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n887), .B1(new_n494), .B2(G128), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n513), .B1(new_n949), .B2(new_n883), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n889), .A2(G164), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n513), .A3(new_n883), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n816), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n850), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n948), .B2(new_n950), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n816), .A3(new_n954), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n848), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n943), .A2(new_n944), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n776), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n943), .A2(new_n775), .A3(new_n944), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n933), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n947), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n947), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n932), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n947), .A2(new_n964), .ZN(new_n968));
  INV_X1    g543(.A(new_n960), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n927), .A2(new_n928), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n659), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n929), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n947), .A2(new_n960), .A3(new_n964), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n967), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT103), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n967), .A2(new_n975), .A3(new_n979), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g557(.A(new_n636), .B1(new_n915), .B2(new_n916), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n538), .B1(new_n527), .B2(new_n528), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n985), .A2(new_n530), .A3(new_n753), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n753), .B1(new_n985), .B2(new_n530), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n602), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n602), .A2(new_n989), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n618), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n992), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(G290), .A3(new_n990), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G305), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n985), .A2(new_n530), .A3(new_n753), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(KEYINPUT105), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n988), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n986), .A2(new_n987), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(KEYINPUT105), .A3(new_n993), .A4(new_n995), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n642), .B(new_n918), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n632), .B(new_n835), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT41), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n632), .A2(G299), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n632), .A2(G299), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n633), .A2(new_n835), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n632), .A2(G299), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(KEYINPUT41), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1008), .B1(new_n1006), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1005), .B(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n983), .B1(new_n1019), .B2(new_n636), .ZN(G295));
  OAI21_X1  g595(.A(new_n983), .B1(new_n1019), .B2(new_n636), .ZN(G331));
  OAI21_X1  g596(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT107), .B1(new_n555), .B2(new_n559), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n914), .A2(new_n917), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n914), .B2(new_n917), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n918), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1022), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n914), .A2(new_n917), .A3(new_n1023), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1026), .A2(new_n1007), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1016), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1035));
  AOI21_X1  g610(.A(G37), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1024), .A2(new_n1025), .A3(new_n1022), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1029), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1012), .B(new_n1015), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1007), .A2(new_n1026), .A3(new_n1031), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1003), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1032), .B1(new_n1040), .B2(KEYINPUT108), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1033), .A2(new_n1046), .A3(new_n1012), .A4(new_n1015), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1035), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n976), .B1(new_n1042), .B2(new_n1003), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT44), .B(new_n1044), .C1(new_n1050), .C2(new_n1037), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT110), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1048), .A2(new_n1049), .A3(KEYINPUT43), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1037), .B1(new_n1036), .B2(new_n1043), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT109), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1040), .A2(KEYINPUT108), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1041), .A3(new_n1047), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1003), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1037), .A3(new_n1036), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT109), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1052), .B1(KEYINPUT44), .B2(new_n1063), .ZN(G397));
  INV_X1    g639(.A(G137), .ZN(new_n1065));
  OAI211_X1 g640(.A(G40), .B(new_n480), .C1(new_n502), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT111), .B1(new_n477), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1069), .B(new_n1066), .C1(new_n469), .C2(new_n476), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1384), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n513), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT45), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n889), .B(new_n892), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1078), .B2(new_n951), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1076), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1080), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT46), .ZN(new_n1082));
  INV_X1    g657(.A(G1996), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n1085), .B(KEYINPUT47), .Z(new_n1086));
  XNOR2_X1  g661(.A(new_n951), .B(G1996), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1076), .B1(new_n1078), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n1088), .B(KEYINPUT112), .Z(new_n1089));
  NOR2_X1   g664(.A1(new_n775), .A2(new_n779), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(new_n1090), .B1(new_n892), .B2(new_n890), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1080), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n776), .A2(new_n778), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1076), .B1(new_n1093), .B2(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT48), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n1080), .A2(G1986), .A3(G290), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT126), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1098), .A2(new_n1096), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1086), .B(new_n1092), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1072), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1075), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1071), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g680(.A(KEYINPUT69), .B(new_n468), .C1(new_n472), .C2(new_n462), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1067), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1069), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n477), .A2(KEYINPUT111), .A3(new_n1067), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n1072), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT45), .B1(new_n513), .B2(new_n1072), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT113), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1105), .A2(new_n765), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1073), .A2(KEYINPUT50), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT50), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n513), .A2(new_n1118), .A3(new_n1072), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1071), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n797), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G8), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(G166), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(G303), .A2(G8), .A3(new_n1124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1123), .A2(G8), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1073), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1126), .B1(new_n1111), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n602), .A2(G1976), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1073), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1131), .B1(new_n602), .B2(G1976), .ZN(new_n1137));
  INV_X1    g712(.A(G1976), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n597), .C1(new_n600), .C2(new_n601), .ZN(new_n1139));
  NOR4_X1   g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .A4(new_n1126), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1981), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n607), .A2(new_n1142), .A3(new_n608), .A4(new_n611), .ZN(new_n1143));
  OAI21_X1  g718(.A(G1981), .B1(new_n751), .B2(new_n752), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT115), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT49), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT49), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1150), .A3(new_n1147), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1133), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT116), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1137), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1133), .A2(new_n1134), .A3(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(G8), .B(new_n1134), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT52), .ZN(new_n1157));
  AND4_X1   g732(.A1(KEYINPUT116), .A2(new_n1152), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1130), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1138), .A3(new_n602), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1143), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1133), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1123), .A2(G8), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1129), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1152), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1123), .A2(G8), .A3(new_n1129), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n878), .B1(new_n1071), .B2(new_n1104), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n513), .A2(new_n1118), .A3(new_n1072), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1118), .B1(new_n513), .B2(new_n1072), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT117), .B(G2084), .Z(new_n1174));
  NAND3_X1  g749(.A1(new_n1111), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1126), .B(G286), .C1(new_n1170), .C2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1167), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1141), .A2(KEYINPUT116), .A3(new_n1152), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1176), .A2(KEYINPUT63), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1183), .A2(new_n1166), .A3(new_n1169), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1163), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1071), .A2(new_n1104), .ZN(new_n1187));
  XNOR2_X1  g762(.A(KEYINPUT56), .B(G2072), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1111), .A2(new_n1173), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT118), .B(G1956), .Z(new_n1190));
  AOI22_X1  g765(.A1(new_n1187), .A2(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT57), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n590), .B1(new_n585), .B2(new_n586), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n554), .B1(new_n575), .B2(new_n576), .ZN(new_n1196));
  INV_X1    g771(.A(new_n589), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1192), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  AND4_X1   g774(.A1(new_n1192), .A2(new_n578), .A3(new_n589), .A4(new_n587), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT119), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT119), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1198), .A2(new_n1192), .A3(new_n587), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT120), .B1(new_n1191), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1136), .A2(new_n892), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(G1348), .B1(new_n1111), .B2(new_n1173), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n633), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1190), .B1(new_n1071), .B2(new_n1120), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1111), .A2(new_n1114), .A3(new_n1188), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT120), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1207), .A2(new_n1211), .A3(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1206), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1111), .A2(new_n1114), .A3(new_n1083), .ZN(new_n1225));
  XNOR2_X1  g800(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(G1341), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1136), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n567), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT59), .ZN(new_n1231));
  OAI211_X1 g806(.A(new_n1231), .B(new_n567), .C1(new_n1225), .C2(new_n1228), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n807), .B1(new_n1071), .B2(new_n1120), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1234), .A2(KEYINPUT60), .A3(new_n1208), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n632), .ZN(new_n1236));
  INV_X1    g811(.A(KEYINPUT60), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1237), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1238));
  NAND4_X1  g813(.A1(new_n1234), .A2(new_n633), .A3(new_n1208), .A4(KEYINPUT60), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1224), .A2(new_n1233), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g816(.A(new_n1217), .ZN(new_n1242));
  OAI21_X1  g817(.A(KEYINPUT61), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1216), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1244));
  NOR3_X1   g819(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1221), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT122), .ZN(new_n1247));
  NOR2_X1   g822(.A1(new_n465), .A2(new_n468), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1247), .B1(new_n1248), .B2(new_n1066), .ZN(new_n1249));
  INV_X1    g824(.A(KEYINPUT53), .ZN(new_n1250));
  NOR2_X1   g825(.A1(new_n1250), .A2(G2078), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NOR3_X1   g827(.A1(new_n1248), .A2(new_n1066), .A3(new_n1247), .ZN(new_n1253));
  NOR2_X1   g828(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI22_X1  g829(.A1(new_n1189), .A2(new_n870), .B1(new_n1114), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g830(.A(G2078), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1256));
  OAI211_X1 g831(.A(G301), .B(new_n1255), .C1(new_n1256), .C2(KEYINPUT53), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1258));
  INV_X1    g833(.A(new_n1251), .ZN(new_n1259));
  OAI22_X1  g834(.A1(new_n1121), .A2(G1961), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NOR3_X1   g835(.A1(new_n1071), .A2(new_n1104), .A3(new_n1102), .ZN(new_n1261));
  AOI21_X1  g836(.A(KEYINPUT113), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1262));
  OAI21_X1  g837(.A(new_n858), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g838(.A(new_n1260), .B1(new_n1263), .B2(new_n1250), .ZN(new_n1264));
  OAI21_X1  g839(.A(new_n1257), .B1(new_n1264), .B2(G301), .ZN(new_n1265));
  INV_X1    g840(.A(KEYINPUT54), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1267));
  NAND2_X1  g842(.A1(new_n1267), .A2(G286), .ZN(new_n1268));
  NAND3_X1  g843(.A1(new_n1170), .A2(G168), .A3(new_n1175), .ZN(new_n1269));
  NAND3_X1  g844(.A1(new_n1268), .A2(G8), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g845(.A1(new_n1270), .A2(KEYINPUT51), .ZN(new_n1271));
  INV_X1    g846(.A(KEYINPUT51), .ZN(new_n1272));
  AND3_X1   g847(.A1(new_n1269), .A2(new_n1272), .A3(G8), .ZN(new_n1273));
  INV_X1    g848(.A(new_n1273), .ZN(new_n1274));
  AOI22_X1  g849(.A1(new_n1265), .A2(new_n1266), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g850(.A(new_n1255), .B1(new_n1256), .B2(KEYINPUT53), .ZN(new_n1276));
  NAND2_X1  g851(.A1(new_n1276), .A2(G171), .ZN(new_n1277));
  INV_X1    g852(.A(new_n1260), .ZN(new_n1278));
  OAI211_X1 g853(.A(new_n1278), .B(G301), .C1(KEYINPUT53), .C2(new_n1256), .ZN(new_n1279));
  NAND3_X1  g854(.A1(new_n1277), .A2(KEYINPUT54), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g855(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1281));
  INV_X1    g856(.A(KEYINPUT124), .ZN(new_n1282));
  NAND4_X1  g857(.A1(new_n1277), .A2(new_n1279), .A3(new_n1282), .A4(KEYINPUT54), .ZN(new_n1283));
  NAND4_X1  g858(.A1(new_n1246), .A2(new_n1275), .A3(new_n1281), .A4(new_n1283), .ZN(new_n1284));
  NAND3_X1  g859(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1285));
  INV_X1    g860(.A(KEYINPUT123), .ZN(new_n1286));
  NAND2_X1  g861(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g862(.A1(new_n1166), .A2(new_n1168), .A3(KEYINPUT123), .A4(new_n1169), .ZN(new_n1288));
  NAND2_X1  g863(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g864(.A(new_n1186), .B1(new_n1284), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g865(.A1(new_n1256), .A2(KEYINPUT53), .ZN(new_n1291));
  OAI21_X1  g866(.A(G171), .B1(new_n1291), .B2(new_n1260), .ZN(new_n1292));
  AOI21_X1  g867(.A(new_n1273), .B1(new_n1270), .B2(KEYINPUT51), .ZN(new_n1293));
  INV_X1    g868(.A(KEYINPUT62), .ZN(new_n1294));
  AOI21_X1  g869(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g870(.A1(new_n1287), .A2(new_n1295), .A3(new_n1288), .ZN(new_n1296));
  INV_X1    g871(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g872(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g873(.A1(new_n1287), .A2(new_n1295), .A3(KEYINPUT125), .A4(new_n1288), .ZN(new_n1299));
  OR2_X1    g874(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1300));
  AND2_X1   g875(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g876(.A(new_n1290), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  AND2_X1   g877(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1303));
  XNOR2_X1  g878(.A(new_n618), .B(G1986), .ZN(new_n1304));
  OAI21_X1  g879(.A(new_n1303), .B1(new_n1080), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g880(.A(new_n1101), .B1(new_n1302), .B2(new_n1305), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g881(.A1(G227), .A2(new_n460), .ZN(new_n1308));
  AOI21_X1  g882(.A(new_n1308), .B1(new_n742), .B2(new_n745), .ZN(new_n1309));
  NAND2_X1  g883(.A1(new_n701), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g884(.A(new_n1310), .B1(new_n978), .B2(new_n980), .ZN(new_n1311));
  AOI21_X1  g885(.A(KEYINPUT127), .B1(new_n1062), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g886(.A(new_n1043), .ZN(new_n1313));
  OAI21_X1  g887(.A(KEYINPUT43), .B1(new_n1313), .B2(new_n1049), .ZN(new_n1314));
  AOI21_X1  g888(.A(new_n1060), .B1(new_n1059), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g889(.A(KEYINPUT109), .B1(new_n1050), .B2(new_n1037), .ZN(new_n1316));
  OAI211_X1 g890(.A(new_n1311), .B(KEYINPUT127), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  INV_X1    g891(.A(new_n1317), .ZN(new_n1318));
  NOR2_X1   g892(.A1(new_n1312), .A2(new_n1318), .ZN(G308));
  OAI21_X1  g893(.A(new_n1311), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1320));
  INV_X1    g894(.A(KEYINPUT127), .ZN(new_n1321));
  NAND2_X1  g895(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g896(.A1(new_n1322), .A2(new_n1317), .ZN(G225));
endmodule


