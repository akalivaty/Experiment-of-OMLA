//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G952), .ZN(new_n187));
  AOI211_X1 g001(.A(G953), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT71), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI211_X1 g008(.A(new_n189), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT21), .B(G898), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n188), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G214), .B1(G237), .B2(G902), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(G210), .B1(G237), .B2(G902), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT0), .B(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(new_n208), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n216), .B2(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n190), .A2(G224), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n218), .B(KEYINPUT92), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT93), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n217), .B(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(G116), .B(G119), .Z(new_n222));
  AND2_X1   g036(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT2), .B(G113), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n223), .B(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT79), .A2(G104), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT79), .A2(G104), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G107), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  INV_X1    g048(.A(G107), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT80), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G107), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G104), .B2(new_n231), .ZN(new_n242));
  OR2_X1    g056(.A1(KEYINPUT79), .A2(G104), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n236), .A3(new_n228), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT80), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n239), .A2(new_n240), .A3(G101), .A4(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(G101), .A3(new_n246), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT81), .A2(G101), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT81), .A2(G101), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n242), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(KEYINPUT4), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT82), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT82), .B1(new_n248), .B2(new_n253), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n227), .B(new_n247), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n243), .A2(new_n235), .A3(new_n228), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n259));
  INV_X1    g073(.A(G101), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(G104), .B2(G107), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n258), .B2(new_n261), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n257), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n264), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n266), .A2(KEYINPUT85), .A3(new_n252), .A4(new_n262), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n222), .A2(new_n224), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n270));
  INV_X1    g084(.A(G119), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G116), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n222), .A2(new_n270), .ZN(new_n275));
  INV_X1    g089(.A(G113), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n269), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n268), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n268), .B2(new_n278), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n256), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT91), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT91), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n256), .B(new_n284), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  XNOR2_X1  g099(.A(G110), .B(G122), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n256), .B(new_n286), .C1(new_n280), .C2(new_n281), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT6), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n286), .B1(new_n282), .B2(KEYINPUT91), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n221), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n265), .A2(new_n267), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n272), .B(KEYINPUT89), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n297));
  OAI21_X1  g111(.A(G113), .B1(new_n222), .B2(new_n297), .ZN(new_n298));
  OAI22_X1  g112(.A1(new_n296), .A2(new_n298), .B1(new_n222), .B2(new_n224), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT94), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  OR3_X1    g114(.A1(new_n295), .A2(KEYINPUT94), .A3(new_n299), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n263), .A2(new_n264), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n278), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n286), .B(KEYINPUT8), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n218), .A2(KEYINPUT7), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n217), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n289), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n189), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n201), .B1(new_n294), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n221), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n292), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n292), .A2(new_n285), .B1(KEYINPUT6), .B2(new_n289), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n307), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n303), .B2(new_n304), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n316), .B2(new_n289), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n200), .A3(new_n317), .ZN(new_n318));
  AOI211_X1 g132(.A(new_n197), .B(new_n199), .C1(new_n310), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT77), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G137), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n321), .A2(KEYINPUT77), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(G125), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n336), .B2(new_n330), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n202), .ZN(new_n338));
  OAI211_X1 g152(.A(G146), .B(new_n332), .C1(new_n336), .C2(new_n330), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n271), .B2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n343), .C1(G119), .C2(new_n213), .ZN(new_n344));
  XNOR2_X1  g158(.A(G119), .B(G128), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT24), .B(G110), .Z(new_n346));
  AOI22_X1  g160(.A1(new_n344), .A2(G110), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n344), .A2(G110), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n339), .C1(G146), .C2(new_n336), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n329), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n325), .A2(new_n348), .A3(new_n350), .A4(new_n328), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n320), .B1(new_n354), .B2(G902), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n352), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n353), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(new_n189), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT78), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(KEYINPUT78), .A3(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(new_n354), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n359), .A2(G902), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT11), .ZN(new_n367));
  INV_X1    g181(.A(G134), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(G137), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT65), .ZN(new_n370));
  INV_X1    g184(.A(G137), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G134), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n367), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G131), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT66), .B1(new_n371), .B2(G134), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT66), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n368), .A3(G137), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n368), .A2(G137), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n377), .A2(new_n379), .B1(new_n380), .B2(KEYINPUT11), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n375), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n376), .B1(new_n375), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n211), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n368), .A2(G137), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n376), .B1(new_n372), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n375), .A2(new_n376), .A3(new_n381), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n215), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(new_n226), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G237), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n194), .A2(G210), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT26), .B(G101), .Z(new_n396));
  OR2_X1    g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n396), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n397), .B2(new_n399), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n384), .A2(new_n226), .A3(KEYINPUT70), .A4(new_n390), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n393), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT73), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n384), .A2(new_n390), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT69), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT64), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n207), .B(new_n410), .C1(new_n208), .C2(new_n209), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n383), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n389), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n390), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n384), .A2(new_n417), .A3(new_n390), .A4(KEYINPUT30), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n408), .A2(new_n416), .A3(new_n227), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n393), .A2(new_n402), .A3(new_n420), .A4(new_n403), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n405), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT31), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n227), .B1(new_n414), .B2(new_n415), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n393), .A2(new_n424), .A3(new_n403), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT28), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n391), .A2(KEYINPUT74), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT74), .B1(new_n391), .B2(new_n427), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n402), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT31), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n405), .A2(new_n434), .A3(new_n419), .A4(new_n421), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n423), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G472), .A2(G902), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n436), .A2(KEYINPUT32), .A3(new_n437), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT75), .B(KEYINPUT32), .Z(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n406), .A2(new_n227), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n393), .A2(new_n403), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT28), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n445), .B2(KEYINPUT28), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n430), .B(new_n443), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n442), .B1(new_n431), .B2(new_n432), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n393), .A2(new_n403), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n419), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n432), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n189), .B(new_n449), .C1(new_n450), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G472), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n366), .B1(new_n441), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  OAI21_X1  g272(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT86), .B(G469), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n194), .A2(G227), .ZN(new_n462));
  XOR2_X1   g276(.A(G110), .B(G140), .Z(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n413), .A2(new_n389), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT10), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n302), .A2(new_n467), .A3(new_n215), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n216), .B1(new_n265), .B2(new_n267), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n467), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n248), .A2(new_n253), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n247), .A2(new_n211), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT83), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT83), .B(new_n476), .C1(new_n254), .C2(new_n255), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n466), .B(new_n470), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n254), .B2(new_n255), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n478), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n466), .B1(new_n485), .B2(new_n470), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT87), .B(new_n464), .C1(new_n481), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n302), .A2(new_n215), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n268), .B2(new_n215), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n465), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT12), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(KEYINPUT12), .A3(new_n465), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n464), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n470), .B1(new_n477), .B2(new_n479), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n465), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n480), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT87), .B1(new_n500), .B2(new_n464), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n189), .B(new_n461), .C1(new_n497), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n480), .A2(new_n495), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n480), .A2(new_n494), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n504), .A2(new_n499), .B1(new_n505), .B2(new_n464), .ZN(new_n506));
  OAI21_X1  g320(.A(G469), .B1(new_n506), .B2(G902), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n460), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT95), .B(G143), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n194), .A2(G214), .A3(new_n394), .A4(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n191), .A2(new_n193), .A3(G214), .A4(new_n394), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n204), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G131), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n513), .A3(new_n376), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT98), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n515), .A2(KEYINPUT98), .A3(new_n516), .A4(new_n517), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n376), .B1(new_n510), .B2(new_n513), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n340), .B1(KEYINPUT17), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G113), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n237), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n510), .B(new_n513), .C1(new_n527), .C2(new_n376), .ZN(new_n528));
  XNOR2_X1  g342(.A(G125), .B(G140), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n202), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n528), .B(new_n530), .C1(new_n515), .C2(new_n527), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n526), .B1(new_n524), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n189), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G475), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n515), .A2(new_n517), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT19), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n336), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n529), .A2(KEYINPUT19), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n339), .B(new_n538), .C1(new_n542), .C2(G146), .ZN(new_n543));
  AOI21_X1  g357(.A(G146), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  INV_X1    g358(.A(new_n339), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT96), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n531), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n526), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(KEYINPUT97), .A3(new_n549), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n532), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT20), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n536), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n213), .A2(G143), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n204), .A2(G128), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT99), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G134), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n563), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n565), .A3(new_n368), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G122), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G116), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n235), .B1(new_n572), .B2(KEYINPUT14), .ZN(new_n573));
  XNOR2_X1  g387(.A(G116), .B(G122), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n563), .B1(new_n577), .B2(new_n565), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n578), .A2(KEYINPUT101), .B1(KEYINPUT13), .B2(new_n566), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n568), .B1(new_n566), .B2(KEYINPUT13), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n368), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n574), .B(new_n235), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n576), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n458), .A2(new_n358), .A3(G953), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n576), .B(new_n587), .C1(new_n583), .C2(new_n585), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT15), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G478), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n560), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n319), .A2(new_n457), .A3(new_n508), .A4(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(new_n251), .Z(G3));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n589), .A2(new_n600), .A3(new_n590), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n589), .B2(new_n590), .ZN(new_n602));
  OAI211_X1 g416(.A(G478), .B(new_n189), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT102), .B(G478), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n591), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n560), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n436), .A2(new_n437), .ZN(new_n609));
  INV_X1    g423(.A(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n436), .B2(new_n189), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n609), .A2(new_n366), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n319), .A2(new_n508), .A3(new_n608), .A4(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  AND2_X1   g429(.A1(new_n508), .A2(new_n612), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n557), .A2(new_n558), .ZN(new_n617));
  INV_X1    g431(.A(new_n534), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n618), .B2(new_n532), .ZN(new_n619));
  INV_X1    g433(.A(G475), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT103), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n535), .A2(new_n622), .A3(G475), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n617), .A2(new_n624), .A3(new_n594), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n616), .A2(new_n319), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  OR2_X1    g442(.A1(new_n609), .A2(new_n611), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n329), .A2(KEYINPUT36), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n630), .A2(KEYINPUT104), .ZN(new_n631));
  INV_X1    g445(.A(new_n351), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(KEYINPUT104), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n635));
  INV_X1    g449(.A(new_n364), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n362), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n637), .A2(new_n638), .A3(new_n360), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n629), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n319), .A3(new_n508), .A4(new_n597), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT105), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT37), .B(G110), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n195), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n188), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n625), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n639), .B1(new_n441), .B2(new_n456), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n199), .B1(new_n310), .B2(new_n318), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n508), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XOR2_X1   g467(.A(new_n647), .B(KEYINPUT39), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n508), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n310), .A2(new_n318), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n436), .A2(KEYINPUT32), .A3(new_n437), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n445), .A2(new_n432), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n422), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n662), .B2(G902), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n660), .B(new_n663), .C1(new_n609), .C2(new_n439), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n560), .A2(new_n595), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n198), .A2(new_n664), .A3(new_n639), .A4(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n656), .A2(new_n657), .A3(new_n659), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  AND3_X1   g482(.A1(new_n559), .A2(new_n606), .A3(new_n648), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n658), .A2(KEYINPUT106), .A3(new_n198), .A4(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n670), .A2(new_n650), .A3(new_n508), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n672));
  INV_X1    g486(.A(new_n651), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n559), .A2(new_n606), .A3(new_n648), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AND2_X1   g491(.A1(new_n502), .A2(new_n459), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n189), .B1(new_n497), .B2(new_n501), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(KEYINPUT107), .A3(G469), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT107), .B1(new_n679), .B2(G469), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(KEYINPUT108), .B(new_n678), .C1(new_n680), .C2(new_n681), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n197), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n651), .A2(new_n687), .A3(new_n608), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n456), .B(new_n660), .C1(new_n609), .C2(new_n439), .ZN(new_n689));
  INV_X1    g503(.A(new_n366), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND4_X1  g509(.A1(new_n658), .A2(new_n625), .A3(new_n687), .A4(new_n198), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n691), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  INV_X1    g513(.A(new_n639), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n689), .A2(new_n597), .A3(new_n687), .A4(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n684), .A2(new_n701), .A3(new_n651), .A4(new_n685), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND3_X1  g517(.A1(new_n651), .A2(new_n687), .A3(new_n665), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n366), .B(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n430), .B1(new_n447), .B2(new_n448), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n432), .B1(KEYINPUT31), .B2(new_n422), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n435), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n432), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n711), .A2(new_n709), .A3(new_n423), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n437), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n436), .A2(new_n189), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT110), .B(G472), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n704), .A2(new_n706), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n684), .A3(new_n685), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND4_X1  g534(.A1(new_n713), .A2(new_n700), .A3(new_n669), .A4(new_n716), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n684), .A2(new_n651), .A3(new_n685), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n310), .A2(new_n318), .A3(new_n198), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n457), .A2(new_n508), .A3(new_n669), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n456), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n436), .A2(new_n437), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT32), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n660), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT112), .A3(new_n660), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n706), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n674), .A2(new_n725), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n726), .A2(new_n508), .A3(new_n737), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n725), .A2(new_n727), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n376), .ZN(G33));
  NAND4_X1  g554(.A1(new_n649), .A2(new_n457), .A3(new_n508), .A4(new_n726), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  NAND2_X1  g556(.A1(new_n560), .A2(new_n606), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT43), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(KEYINPUT43), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n629), .A3(new_n700), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(G469), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n505), .A2(new_n464), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n503), .B2(new_n486), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n506), .A2(KEYINPUT45), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n753), .A2(new_n754), .B1(G469), .B2(G902), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n502), .B1(new_n755), .B2(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n459), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n310), .A2(new_n318), .A3(new_n198), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n746), .B2(new_n747), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n748), .A2(new_n759), .A3(new_n654), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT113), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n689), .A2(new_n760), .A3(new_n690), .A4(new_n674), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n766), .B(new_n767), .C1(new_n758), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  AND2_X1   g584(.A1(new_n686), .A2(new_n726), .ZN(new_n771));
  INV_X1    g585(.A(new_n188), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n664), .A2(new_n366), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n560), .A3(new_n607), .A4(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n713), .A2(new_n716), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n744), .A2(new_n188), .A3(new_n745), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n771), .A2(new_n700), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n366), .B(KEYINPUT111), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n776), .A2(new_n779), .A3(new_n775), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n659), .A2(new_n198), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n686), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT50), .Z(new_n783));
  AND2_X1   g597(.A1(new_n780), .A2(new_n726), .ZN(new_n784));
  INV_X1    g598(.A(new_n766), .ZN(new_n785));
  INV_X1    g599(.A(new_n768), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n759), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n680), .A2(new_n681), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n460), .A3(new_n502), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n784), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n778), .A2(new_n783), .A3(KEYINPUT51), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n771), .A2(new_n608), .A3(new_n773), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n780), .A2(new_n686), .A3(new_n651), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(G952), .A3(new_n190), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n771), .A2(new_n776), .ZN(new_n796));
  INV_X1    g610(.A(new_n736), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n796), .A2(KEYINPUT48), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT48), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n789), .B(KEYINPUT116), .Z(new_n801));
  OAI21_X1  g615(.A(new_n784), .B1(new_n787), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n778), .A2(new_n783), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n792), .B(new_n800), .C1(new_n803), .C2(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n502), .A2(new_n507), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n637), .A2(new_n638), .A3(new_n360), .A4(new_n647), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n664), .A3(new_n459), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n651), .A2(new_n665), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n671), .B2(new_n675), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n723), .A3(new_n652), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n594), .B(new_n536), .C1(new_n558), .C2(new_n557), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n658), .A2(new_n687), .A3(new_n198), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n651), .A2(new_n818), .A3(new_n687), .A4(new_n815), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n616), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n598), .A3(new_n613), .A4(new_n641), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n617), .A2(new_n624), .A3(new_n595), .A4(new_n648), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n689), .A2(new_n822), .A3(new_n700), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n721), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n805), .A2(new_n459), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n760), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n741), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n821), .A2(new_n739), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n810), .A2(new_n723), .A3(new_n830), .A4(new_n652), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n684), .B(new_n685), .C1(new_n692), .C2(new_n697), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(new_n702), .A3(new_n719), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n813), .A2(new_n829), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n829), .A3(new_n831), .A4(new_n833), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT54), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n835), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n832), .A2(new_n719), .A3(new_n702), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n727), .A2(new_n725), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n736), .A2(new_n738), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n691), .A2(new_n825), .A3(new_n760), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n846), .A2(new_n649), .B1(new_n824), .B2(new_n826), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n842), .A2(new_n848), .A3(new_n821), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT53), .A3(new_n831), .A4(new_n813), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n841), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n804), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n788), .A2(new_n502), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT49), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n779), .A2(new_n459), .A3(new_n198), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n659), .A2(new_n858), .A3(new_n664), .A4(new_n743), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(KEYINPUT49), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n854), .A2(new_n855), .B1(new_n857), .B2(new_n861), .ZN(G75));
  INV_X1    g676(.A(new_n194), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n187), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT118), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n841), .A2(new_n850), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(G902), .ZN(new_n869));
  INV_X1    g683(.A(G210), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n291), .A2(new_n293), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT117), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n221), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n875), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n867), .B(new_n877), .C1(new_n869), .C2(new_n870), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n866), .B1(new_n876), .B2(new_n878), .ZN(G51));
  INV_X1    g693(.A(new_n852), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n851), .B1(new_n841), .B2(new_n850), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(G469), .A2(G902), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT57), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n882), .A2(new_n884), .B1(new_n501), .B2(new_n497), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n189), .B1(new_n841), .B2(new_n850), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n753), .A2(new_n754), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(KEYINPUT119), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT119), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n866), .B1(new_n885), .B2(new_n891), .ZN(G54));
  AND4_X1   g706(.A1(KEYINPUT58), .A2(new_n868), .A3(G475), .A4(G902), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n865), .B1(new_n893), .B2(new_n554), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .A4(new_n554), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT120), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n895), .A2(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G60));
  OR2_X1    g712(.A1(new_n601), .A2(new_n602), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT59), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n853), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n865), .B1(new_n882), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n868), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n866), .B1(new_n909), .B2(new_n354), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n841), .B2(new_n850), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n634), .A2(new_n635), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n910), .A2(KEYINPUT121), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n865), .B1(new_n912), .B2(new_n363), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n913), .B(new_n907), .C1(new_n841), .C2(new_n850), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n916), .A2(new_n921), .ZN(G66));
  INV_X1    g736(.A(G224), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n196), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n842), .A2(new_n821), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n863), .ZN(new_n926));
  INV_X1    g740(.A(G898), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n873), .B1(new_n927), .B2(new_n863), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n926), .B(new_n928), .Z(G69));
  INV_X1    g743(.A(G227), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n863), .B1(new_n930), .B2(new_n645), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT124), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n769), .A2(new_n762), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n723), .A2(new_n652), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n676), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n759), .A2(new_n654), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n736), .A2(new_n651), .A3(new_n665), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n845), .B(new_n741), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n934), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n194), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n408), .A2(new_n416), .A3(new_n418), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT122), .Z(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(new_n542), .Z(new_n944));
  OAI211_X1 g758(.A(new_n941), .B(new_n944), .C1(new_n645), .C2(new_n194), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n457), .B(new_n726), .C1(new_n608), .C2(new_n815), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(new_n655), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n769), .A2(new_n762), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n935), .A2(new_n667), .A3(new_n676), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n944), .B1(new_n954), .B2(new_n194), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n945), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(KEYINPUT123), .B(new_n944), .C1(new_n954), .C2(new_n194), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n933), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n950), .A2(new_n951), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n950), .A2(new_n951), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n948), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n863), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT123), .B1(new_n963), .B2(new_n944), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n955), .A2(new_n956), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n965), .A3(new_n932), .A4(new_n945), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n959), .A2(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n962), .B2(new_n925), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n452), .B(KEYINPUT125), .Z(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n432), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n453), .B2(new_n422), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT126), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n839), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n970), .B1(new_n940), .B2(new_n925), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n972), .A2(new_n432), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n865), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n973), .A2(new_n976), .A3(new_n979), .ZN(G57));
endmodule


