//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT29), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT79), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n207), .A2(new_n208), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n209), .A2(new_n212), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n216), .A2(new_n218), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(new_n220), .A3(new_n212), .A4(new_n209), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  AND2_X1   g024(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n231), .B(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT67), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n226), .A2(new_n227), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT28), .A3(new_n225), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n229), .A2(new_n238), .A3(new_n230), .A4(new_n232), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n215), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n213), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n242), .B1(new_n210), .B2(new_n241), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n206), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(KEYINPUT69), .B(new_n206), .C1(new_n245), .C2(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI221_X4 g050(.A(new_n205), .B1(new_n222), .B2(new_n224), .C1(new_n240), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(new_n251), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n222), .A2(new_n224), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT79), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n204), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n262), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n240), .A2(new_n251), .B1(new_n222), .B2(new_n224), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n203), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n256), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n252), .A2(new_n255), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n254), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n270), .A2(new_n203), .B1(new_n204), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT80), .B(new_n269), .C1(new_n272), .C2(new_n266), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n274), .A3(new_n266), .A4(new_n268), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n273), .A2(new_n275), .A3(new_n279), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n271), .A2(new_n205), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n267), .A2(KEYINPUT79), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n203), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n204), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n274), .B1(new_n289), .B2(new_n265), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(new_n269), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n291), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(G148gat), .ZN(new_n295));
  INV_X1    g094(.A(G148gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(G141gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G155gat), .B2(G162gat), .ZN(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT81), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n298), .A2(new_n299), .A3(new_n301), .A4(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT71), .B(KEYINPUT1), .ZN(new_n307));
  INV_X1    g106(.A(G113gat), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n309), .A2(G113gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n306), .B(new_n307), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n308), .A2(G120gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n306), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n293), .A2(new_n302), .A3(new_n303), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n299), .ZN(new_n322));
  OR2_X1    g121(.A1(KEYINPUT82), .A2(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(KEYINPUT82), .A2(G141gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n296), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(new_n325), .B2(new_n295), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n305), .A2(new_n315), .A3(new_n320), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT4), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n296), .A2(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n294), .A2(G148gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT2), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n301), .ZN(new_n332));
  INV_X1    g131(.A(new_n299), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n324), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT82), .A2(G141gat), .ZN(new_n336));
  OAI21_X1  g135(.A(G148gat), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n337), .A2(new_n329), .B1(new_n299), .B2(new_n321), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n306), .A2(new_n307), .ZN(new_n341));
  INV_X1    g140(.A(new_n314), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT70), .B(G120gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(new_n308), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n341), .A2(new_n344), .B1(new_n318), .B2(new_n319), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n346), .A3(KEYINPUT85), .ZN(new_n347));
  OR3_X1    g146(.A1(new_n327), .A2(KEYINPUT85), .A3(KEYINPUT4), .ZN(new_n348));
  INV_X1    g147(.A(new_n345), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n334), .B2(new_n338), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n305), .A2(new_n351), .A3(new_n326), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT83), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n305), .A2(new_n326), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n327), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n357), .B(KEYINPUT39), .C1(new_n356), .C2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G1gat), .B(G29gat), .Z(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(G85gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G57gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n361), .B(new_n365), .C1(KEYINPUT39), .C2(new_n357), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT40), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(new_n360), .B2(new_n356), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n327), .B2(KEYINPUT4), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n339), .A2(KEYINPUT84), .A3(new_n345), .A4(new_n340), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n372), .A2(new_n373), .A3(new_n328), .ZN(new_n374));
  INV_X1    g173(.A(new_n356), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n378), .A2(new_n369), .A3(new_n348), .A4(new_n347), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n365), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n368), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n367), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n283), .A2(new_n292), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT90), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n377), .A2(new_n365), .A3(new_n379), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n382), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT91), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n365), .B(new_n389), .C1(new_n377), .C2(new_n379), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n380), .B2(new_n381), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n393), .B1(new_n394), .B2(new_n390), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n395), .B2(KEYINPUT91), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT37), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n280), .B1(new_n276), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n256), .A2(new_n265), .A3(new_n268), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n272), .B2(new_n265), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n397), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(KEYINPUT38), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n396), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n279), .B1(new_n291), .B2(KEYINPUT37), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n273), .A2(KEYINPUT37), .A3(new_n275), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT38), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n406), .A3(new_n281), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n262), .A2(new_n264), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n263), .B1(new_n261), .B2(new_n257), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n339), .B1(new_n351), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n265), .B1(new_n408), .B2(new_n352), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT87), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT87), .B(new_n415), .C1(new_n412), .C2(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n421), .A3(new_n418), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT88), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n421), .B1(new_n417), .B2(new_n418), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT89), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n422), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n431), .B2(new_n427), .ZN(new_n432));
  INV_X1    g231(.A(new_n426), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n420), .B2(KEYINPUT88), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n422), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n430), .A2(new_n436), .B1(new_n437), .B2(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n283), .A2(new_n292), .A3(new_n385), .A4(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n387), .A2(new_n407), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n253), .A2(new_n345), .A3(new_n254), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT72), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n271), .A2(new_n349), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n345), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT73), .B(KEYINPUT33), .Z(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  INV_X1    g255(.A(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT74), .B(G71gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT32), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n449), .B2(new_n451), .ZN(new_n464));
  INV_X1    g263(.A(new_n454), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n449), .B2(new_n451), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n466), .B2(new_n460), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n446), .A2(new_n447), .A3(new_n450), .A4(new_n448), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n450), .B2(KEYINPUT76), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT77), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n468), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n462), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT78), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n462), .A2(new_n476), .A3(new_n467), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT75), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n464), .A2(new_n466), .A3(new_n460), .ZN(new_n480));
  AOI221_X4 g279(.A(new_n463), .B1(new_n461), .B2(new_n465), .C1(new_n449), .C2(new_n451), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n462), .A2(KEYINPUT75), .A3(new_n467), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n443), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n473), .B1(new_n462), .B2(new_n467), .ZN(new_n487));
  AOI211_X1 g286(.A(KEYINPUT36), .B(new_n487), .C1(new_n475), .C2(new_n477), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n283), .A2(new_n292), .ZN(new_n490));
  INV_X1    g289(.A(new_n395), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n439), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n442), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n439), .A3(new_n485), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n282), .A2(KEYINPUT30), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n279), .B1(new_n273), .B2(new_n275), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n291), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n487), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT92), .B1(new_n478), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504));
  AOI211_X1 g303(.A(new_n504), .B(new_n487), .C1(new_n475), .C2(new_n477), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n490), .A2(new_n507), .A3(new_n439), .A4(new_n396), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n501), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G8gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT97), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518));
  AOI21_X1  g317(.A(G8gat), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n513), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G50gat), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n523), .A2(G43gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(G43gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT15), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT95), .B(G43gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n523), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT15), .B1(new_n528), .B2(new_n524), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  OAI22_X1  g333(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n526), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n526), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT17), .B1(new_n539), .B2(KEYINPUT96), .ZN(new_n540));
  AND4_X1   g339(.A1(KEYINPUT96), .A2(new_n536), .A3(KEYINPUT17), .A4(new_n537), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n522), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n517), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n539), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT99), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT18), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n522), .A2(new_n538), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n544), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n545), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(KEYINPUT99), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G113gat), .B(G141gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT94), .ZN(new_n557));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n562), .A3(new_n552), .A4(new_n554), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT7), .ZN(new_n568));
  INV_X1    g367(.A(G106gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT8), .B1(new_n457), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT101), .B(G85gat), .Z(new_n571));
  OAI211_X1 g370(.A(new_n568), .B(new_n570), .C1(G92gat), .C2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G57gat), .B(G64gat), .Z(new_n575));
  INV_X1    g374(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n573), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n572), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G230gat), .ZN(new_n594));
  INV_X1    g393(.A(G233gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n585), .A2(new_n589), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n596), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT100), .Z(new_n611));
  AOI21_X1  g410(.A(new_n543), .B1(KEYINPUT21), .B2(new_n588), .ZN(new_n612));
  INV_X1    g411(.A(G183gat), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n616), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n623));
  INV_X1    g422(.A(new_n611), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n584), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n259), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n620), .A2(new_n625), .A3(new_n631), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n574), .B1(new_n540), .B2(new_n541), .ZN(new_n639));
  NAND3_X1  g438(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n639), .B(new_n640), .C1(new_n538), .C2(new_n574), .ZN(new_n641));
  XOR2_X1   g440(.A(G190gat), .B(G218gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n638), .B1(new_n644), .B2(KEYINPUT102), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n643), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g449(.A1(new_n510), .A2(new_n566), .A3(new_n609), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n395), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(G1gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  INV_X1    g453(.A(new_n490), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  AOI21_X1  g456(.A(KEYINPUT42), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT104), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(KEYINPUT42), .A3(new_n657), .ZN(new_n660));
  INV_X1    g459(.A(G8gat), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n659), .B(new_n660), .C1(new_n661), .C2(new_n656), .ZN(G1325gat));
  INV_X1    g461(.A(new_n506), .ZN(new_n663));
  AOI21_X1  g462(.A(G15gat), .B1(new_n651), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n489), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n651), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(G15gat), .B2(new_n666), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n438), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n649), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n494), .B2(new_n509), .ZN(new_n672));
  INV_X1    g471(.A(new_n635), .ZN(new_n673));
  INV_X1    g472(.A(new_n566), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n673), .A2(new_n674), .A3(new_n608), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n533), .A3(new_n395), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n675), .B(KEYINPUT105), .Z(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n510), .A2(new_n649), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n672), .A2(KEYINPUT108), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n672), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n492), .A2(new_n486), .A3(new_n488), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT35), .B(new_n438), .C1(new_n283), .C2(new_n292), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n691), .B(new_n396), .C1(new_n503), .C2(new_n505), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n690), .A2(new_n442), .B1(new_n692), .B2(new_n501), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n693), .C2(new_n671), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n679), .B1(new_n686), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(new_n395), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n678), .B1(new_n697), .B2(new_n533), .ZN(G1328gat));
  NAND3_X1  g497(.A1(new_n676), .A2(new_n534), .A3(new_n655), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT46), .Z(new_n700));
  AND2_X1   g499(.A1(new_n696), .A2(new_n655), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n534), .ZN(G1329gat));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  INV_X1    g502(.A(new_n527), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n676), .A2(new_n663), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n704), .B1(new_n696), .B2(new_n665), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n696), .A2(new_n665), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT47), .B(new_n706), .C1(new_n710), .C2(new_n704), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(G1330gat));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  AOI211_X1 g512(.A(new_n439), .B(new_n679), .C1(new_n686), .C2(new_n695), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n523), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n676), .A2(new_n523), .A3(new_n438), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n714), .B2(new_n523), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI221_X1 g518(.A(new_n716), .B1(new_n713), .B2(KEYINPUT48), .C1(new_n714), .C2(new_n523), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1331gat));
  NAND3_X1  g520(.A1(new_n650), .A2(new_n674), .A3(new_n608), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT111), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n510), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n395), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g526(.A1(new_n724), .A2(KEYINPUT112), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(KEYINPUT112), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n490), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n489), .B1(new_n728), .B2(new_n729), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(new_n577), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n725), .A2(new_n577), .A3(new_n663), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(new_n738), .C1(new_n736), .C2(new_n577), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(G1334gat));
  AOI21_X1  g541(.A(new_n439), .B1(new_n728), .B2(new_n729), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT113), .B(G78gat), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n673), .A2(new_n566), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n686), .B2(new_n695), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n395), .A3(new_n608), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT114), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n748), .A2(new_n751), .A3(new_n395), .A4(new_n608), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n571), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n672), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT51), .B1(new_n754), .B2(new_n747), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n755), .A2(new_n608), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n491), .A2(new_n571), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(G1336gat));
  NAND4_X1  g559(.A1(new_n755), .A2(new_n655), .A3(new_n608), .A4(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(G92gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n748), .A2(G92gat), .A3(new_n608), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n490), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(KEYINPUT52), .B(new_n763), .C1(new_n764), .C2(new_n490), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n757), .A2(new_n457), .A3(new_n663), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n748), .A2(new_n665), .A3(new_n608), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n457), .ZN(G1338gat));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n438), .A3(new_n608), .A4(new_n756), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n569), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n748), .A2(G106gat), .A3(new_n608), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n439), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(KEYINPUT53), .B(new_n774), .C1(new_n775), .C2(new_n439), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n596), .B1(new_n591), .B2(new_n592), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n606), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT54), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n782), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n781), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n784), .B(KEYINPUT55), .C1(new_n782), .C2(new_n787), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n607), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT115), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n789), .A2(new_n607), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n792), .A2(new_n794), .B1(new_n564), .B2(new_n565), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n550), .A2(new_n551), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n545), .B1(new_n542), .B2(new_n544), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n561), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n565), .A2(new_n608), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n671), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n794), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n565), .A2(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n649), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n673), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n635), .A2(new_n649), .A3(new_n566), .A4(new_n608), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n806), .B2(new_n438), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n439), .C1(new_n804), .C2(new_n805), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n506), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n655), .A2(new_n491), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n674), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n806), .A2(new_n438), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n478), .A2(new_n485), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n811), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n308), .A3(new_n566), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n819), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n812), .B2(new_n609), .ZN(new_n821));
  INV_X1    g620(.A(new_n343), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n822), .A3(new_n608), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1341gat));
  AOI21_X1  g623(.A(G127gat), .B1(new_n818), .B2(new_n673), .ZN(new_n825));
  INV_X1    g624(.A(new_n812), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n673), .A2(G127gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(G1342gat));
  INV_X1    g627(.A(G134gat), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n829), .A3(new_n815), .A4(new_n811), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n671), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT56), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n649), .A3(new_n811), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT117), .B1(new_n833), .B2(G134gat), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n833), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n832), .B(KEYINPUT118), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n335), .A2(new_n336), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n799), .A2(KEYINPUT119), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n799), .A2(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n674), .A2(new_n791), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n671), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n673), .B1(new_n846), .B2(new_n803), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n438), .C1(new_n847), .C2(new_n805), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n650), .A2(new_n674), .A3(new_n609), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n842), .B(new_n843), .C1(new_n674), .C2(new_n791), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n649), .A2(new_n802), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n851), .A2(new_n671), .B1(new_n801), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n853), .B2(new_n673), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT57), .A4(new_n438), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n806), .B2(new_n439), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n849), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n665), .A2(new_n817), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n841), .B1(new_n861), .B2(new_n674), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n806), .A2(new_n439), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n860), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n294), .A3(new_n566), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n862), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1344gat));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n296), .A3(new_n608), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n861), .B2(new_n609), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n296), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n852), .A2(new_n607), .A3(new_n790), .A4(new_n789), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n673), .B1(new_n846), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n857), .B(new_n438), .C1(new_n877), .C2(new_n805), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n806), .B2(new_n439), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n608), .A3(new_n860), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n873), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n872), .B1(new_n875), .B2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(new_n302), .B1(new_n864), .B2(new_n635), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n859), .A2(G155gat), .A3(new_n860), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n635), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT121), .ZN(G1346gat));
  AOI21_X1  g686(.A(G162gat), .B1(new_n865), .B2(new_n649), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n861), .A2(new_n671), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n490), .A2(new_n395), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n816), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G169gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n566), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n799), .B1(new_n801), .B2(new_n566), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n803), .B1(new_n896), .B2(new_n649), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n635), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n850), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n808), .B1(new_n899), .B2(new_n439), .ZN(new_n900));
  INV_X1    g699(.A(new_n809), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n663), .B(new_n891), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n807), .A2(new_n809), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n663), .A4(new_n891), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n904), .A2(new_n566), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n895), .B1(new_n907), .B2(new_n894), .ZN(G1348gat));
  AOI21_X1  g707(.A(G176gat), .B1(new_n893), .B2(new_n608), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n904), .A2(new_n608), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(G176gat), .ZN(G1349gat));
  OR2_X1    g710(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n904), .A2(new_n673), .A3(new_n906), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G183gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n816), .A2(new_n235), .A3(new_n635), .A4(new_n892), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n912), .A2(new_n914), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n913), .B2(G183gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n912), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n920), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n893), .A2(new_n225), .A3(new_n649), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n649), .A3(new_n906), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(G190gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n923), .B2(G190gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n665), .A2(new_n892), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n880), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n674), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n490), .A2(new_n439), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n489), .A2(KEYINPUT124), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT124), .B1(new_n489), .B2(new_n931), .ZN(new_n933));
  NOR4_X1   g732(.A1(new_n806), .A2(new_n932), .A3(new_n933), .A4(new_n395), .ZN(new_n934));
  INV_X1    g733(.A(G197gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n935), .A3(new_n566), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n930), .A2(new_n936), .ZN(G1352gat));
  INV_X1    g736(.A(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n938), .A3(new_n608), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT126), .B1(new_n943), .B2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n880), .A2(new_n608), .A3(new_n928), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G204gat), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n941), .A2(new_n948), .A3(new_n949), .A4(new_n942), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n944), .A2(new_n945), .A3(new_n947), .A4(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n259), .A3(new_n673), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n880), .A2(new_n673), .A3(new_n928), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  AOI21_X1  g755(.A(G218gat), .B1(new_n934), .B2(new_n649), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n929), .A2(new_n671), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(G218gat), .ZN(G1355gat));
endmodule


