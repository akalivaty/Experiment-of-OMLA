//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT73), .B1(new_n204), .B2(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(G141gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(G141gat), .C2(new_n207), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n213), .B2(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n204), .A2(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n207), .A2(G141gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n213), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT71), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(KEYINPUT71), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G211gat), .B(G218gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n228), .A3(new_n225), .A4(new_n226), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT29), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n222), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n214), .A2(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT77), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n231), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI211_X1 g041(.A(KEYINPUT77), .B(KEYINPUT29), .C1(new_n234), .C2(new_n235), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n203), .B(new_n233), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n233), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n202), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT78), .B(G22gat), .Z(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT79), .ZN(new_n250));
  XOR2_X1   g049(.A(G78gat), .B(G106gat), .Z(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT31), .B(G50gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n254), .B1(new_n236), .B2(new_n237), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n255), .A2(new_n243), .A3(new_n240), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n233), .A2(new_n203), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n247), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n253), .B1(new_n258), .B2(G22gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n247), .A3(new_n260), .A4(new_n248), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n250), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n249), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n248), .B1(new_n244), .B2(new_n247), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n253), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(KEYINPUT23), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G169gat), .ZN(new_n272));
  INV_X1    g071(.A(G176gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n273), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT25), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT24), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n281), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n294), .A3(new_n275), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n267), .A2(KEYINPUT23), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n275), .A2(new_n280), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n286), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n274), .B1(KEYINPUT26), .B2(new_n278), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT26), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n269), .A2(new_n306), .A3(new_n270), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n308), .A2(new_n282), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT67), .B(G183gat), .ZN(new_n310));
  AOI21_X1  g109(.A(G190gat), .B1(new_n310), .B2(KEYINPUT27), .ZN(new_n311));
  OR2_X1    g110(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n312));
  NAND2_X1  g111(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(G183gat), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT28), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT27), .B(G183gat), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n316), .A2(new_n317), .A3(G190gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n309), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G226gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n320), .B2(new_n237), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n241), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n315), .ZN(new_n331));
  INV_X1    g130(.A(new_n318), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n333), .A2(new_n309), .B1(new_n296), .B2(new_n303), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n334), .A2(KEYINPUT29), .B1(new_n321), .B2(new_n322), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(new_n240), .A3(new_n324), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(KEYINPUT1), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G113gat), .B(G120gat), .Z(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n234), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n348), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n222), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n341), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT75), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n234), .B(new_n351), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(KEYINPUT5), .C1(new_n357), .C2(new_n341), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT74), .B1(new_n234), .B2(new_n235), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n222), .A2(new_n360), .A3(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n349), .B1(new_n235), .B2(new_n234), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n341), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT69), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT69), .B1(new_n344), .B2(new_n348), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n234), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(KEYINPUT4), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n355), .B(new_n358), .C1(new_n365), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n234), .C1(new_n367), .C2(new_n368), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n372), .A2(new_n374), .B1(new_n362), .B2(new_n363), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT5), .B1(G225gat), .B2(G233gat), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT76), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n372), .ZN(new_n378));
  AND4_X1   g177(.A1(KEYINPUT76), .A2(new_n378), .A3(new_n364), .A4(new_n376), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n371), .B(new_n384), .C1(new_n377), .C2(new_n379), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n340), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n330), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n325), .A2(new_n326), .A3(new_n241), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n240), .B1(new_n335), .B2(new_n324), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n327), .A2(new_n336), .A3(KEYINPUT30), .A4(new_n330), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n266), .B1(new_n391), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT36), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n367), .A2(new_n368), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n301), .B1(new_n298), .B2(new_n299), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n294), .B1(new_n271), .B2(new_n275), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n292), .A2(new_n286), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(new_n281), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n408), .B2(new_n295), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n308), .A2(new_n282), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n331), .B2(new_n332), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G227gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n322), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n304), .A2(new_n319), .A3(new_n403), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G15gat), .B(G43gat), .Z(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n416), .B(KEYINPUT32), .C1(new_n418), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT70), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n415), .ZN(new_n429));
  INV_X1    g228(.A(new_n414), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT34), .B(new_n414), .C1(new_n412), .C2(new_n415), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n433), .A2(new_n423), .A3(new_n425), .ZN(new_n434));
  INV_X1    g233(.A(new_n431), .ZN(new_n435));
  INV_X1    g234(.A(new_n432), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n423), .A2(new_n425), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n427), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(KEYINPUT70), .A3(new_n433), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n402), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n437), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n423), .A3(new_n425), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT36), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n401), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT37), .B1(new_n393), .B2(new_n394), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n327), .A2(new_n447), .A3(new_n336), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n392), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT83), .B(KEYINPUT38), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n446), .A2(new_n392), .A3(new_n448), .A4(new_n450), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n389), .A2(new_n390), .A3(new_n337), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n395), .A2(new_n397), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n339), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n395), .A2(new_n397), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT80), .B1(new_n340), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n341), .B1(new_n378), .B2(new_n364), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n385), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n357), .B2(new_n341), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n375), .B2(new_n341), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT82), .A4(KEYINPUT40), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT81), .B(KEYINPUT40), .Z(new_n474));
  AOI22_X1  g273(.A1(new_n385), .A2(new_n380), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n456), .A2(new_n477), .A3(new_n266), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n391), .A2(new_n400), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n438), .A2(new_n266), .A3(new_n439), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT35), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n389), .A2(new_n390), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n434), .A2(new_n437), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT35), .B1(new_n262), .B2(new_n265), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(new_n462), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n445), .A2(new_n478), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G197gat), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT11), .B(G169gat), .Z(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT12), .ZN(new_n492));
  INV_X1    g291(.A(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT16), .ZN(new_n494));
  INV_X1    g293(.A(G15gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(G22gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G15gat), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(G1gat), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g299(.A(G8gat), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n502), .B(new_n503), .C1(G1gat), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G43gat), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G50gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  AND2_X1   g312(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n512), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n509), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n510), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n516), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n526), .B2(new_n512), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT17), .B1(new_n527), .B2(KEYINPUT86), .ZN(new_n528));
  INV_X1    g327(.A(new_n512), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n524), .B2(new_n525), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NOR4_X1   g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n519), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n507), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n526), .A2(new_n512), .ZN(new_n536));
  INV_X1    g335(.A(new_n519), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n536), .A2(new_n537), .A3(new_n506), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n535), .A4(new_n539), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n535), .B(KEYINPUT13), .Z(new_n544));
  AOI21_X1  g343(.A(new_n506), .B1(new_n536), .B2(new_n537), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT87), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT87), .B(new_n544), .C1(new_n538), .C2(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND4_X1   g349(.A1(new_n492), .A2(new_n542), .A3(new_n543), .A4(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n540), .A2(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n492), .B1(new_n552), .B2(new_n543), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n528), .A2(new_n533), .ZN(new_n555));
  AND2_X1   g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  AND2_X1   g355(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(KEYINPUT93), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT7), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT8), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(G99gat), .B2(G106gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G99gat), .ZN(new_n575));
  INV_X1    g374(.A(G106gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT8), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n573), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT94), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n568), .A2(new_n569), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n569), .B1(new_n568), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n555), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n527), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT41), .ZN(new_n586));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n584), .A2(new_n588), .B1(KEYINPUT95), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n586), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT90), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(KEYINPUT95), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n593), .A2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G230gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n322), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G57gat), .B(G64gat), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(G71gat), .A2(G78gat), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n604), .A2(new_n605), .B1(KEYINPUT88), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G71gat), .B(G78gat), .Z(new_n608));
  AND2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n581), .B2(new_n582), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n563), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n567), .B1(new_n617), .B2(KEYINPUT93), .ZN(new_n618));
  INV_X1    g417(.A(new_n562), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n580), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n569), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n607), .B(new_n608), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n568), .A2(new_n569), .A3(new_n580), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n603), .B1(new_n612), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n612), .A2(new_n625), .A3(new_n631), .A4(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(new_n625), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n630), .A2(new_n632), .B1(new_n633), .B2(KEYINPUT10), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n627), .B1(new_n634), .B2(new_n602), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT21), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n611), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G127gat), .B(G155gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n507), .B1(new_n611), .B2(new_n645), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT89), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n650), .B(new_n656), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n600), .A2(new_n644), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT98), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n600), .A2(new_n644), .A3(new_n660), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n487), .A2(new_n554), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n482), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n462), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT99), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(G8gat), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND4_X1  g470(.A1(new_n663), .A2(KEYINPUT42), .A3(new_n462), .A4(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(new_n671), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n673), .B(KEYINPUT100), .C1(new_n675), .C2(KEYINPUT42), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT42), .B1(new_n674), .B2(new_n671), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n670), .A2(new_n672), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(G1325gat));
  INV_X1    g480(.A(new_n663), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n440), .A2(new_n444), .ZN(new_n683));
  OAI21_X1  g482(.A(G15gat), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n663), .A2(new_n495), .A3(new_n483), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1326gat));
  INV_X1    g485(.A(new_n266), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n487), .B2(new_n600), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n593), .B(new_n597), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n479), .A2(new_n687), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n438), .A2(new_n439), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT36), .ZN(new_n696));
  INV_X1    g495(.A(new_n444), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n266), .B1(new_n454), .B2(new_n455), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n473), .A2(new_n475), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n461), .B2(new_n459), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n481), .A2(new_n486), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n693), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n692), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n657), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n551), .B2(new_n553), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n542), .A2(new_n543), .A3(new_n550), .ZN(new_n710));
  INV_X1    g509(.A(new_n492), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n552), .A2(new_n492), .A3(new_n543), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT101), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n707), .A2(new_n644), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n482), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n693), .A2(new_n707), .A3(new_n644), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n487), .A2(new_n554), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n517), .A3(new_n664), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1328gat));
  INV_X1    g522(.A(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(new_n462), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n724), .A2(G36gat), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(KEYINPUT102), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n717), .B2(new_n725), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G36gat), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n730), .A3(new_n725), .ZN(new_n733));
  OAI221_X1 g532(.A(new_n728), .B1(new_n726), .B2(new_n729), .C1(new_n732), .C2(new_n733), .ZN(G1329gat));
  NOR3_X1   g533(.A1(new_n724), .A2(G43gat), .A3(new_n443), .ZN(new_n735));
  INV_X1    g534(.A(new_n683), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n706), .A2(new_n736), .A3(new_n716), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g538(.A1(new_n692), .A2(new_n705), .A3(new_n687), .A4(new_n716), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n266), .A2(G50gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n720), .A2(new_n743), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n741), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n747), .B(new_n749), .ZN(G1331gat));
  INV_X1    g549(.A(new_n644), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n600), .A2(new_n751), .A3(new_n657), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n487), .A2(new_n715), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n664), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g554(.A(new_n753), .B(KEYINPUT106), .Z(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n725), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n756), .B2(new_n683), .ZN(new_n762));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n753), .A2(KEYINPUT107), .A3(new_n483), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n753), .B2(new_n483), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1334gat));
  NOR2_X1   g568(.A1(new_n756), .A2(new_n266), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(G78gat), .Z(G1335gat));
  INV_X1    g570(.A(new_n487), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n715), .A2(new_n657), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n693), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n693), .A4(new_n773), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n644), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(G85gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n664), .ZN(new_n780));
  INV_X1    g579(.A(new_n773), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n644), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n692), .A2(new_n705), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT108), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n692), .A2(new_n705), .A3(new_n785), .A4(new_n782), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n784), .A2(new_n664), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n780), .B1(new_n787), .B2(new_n779), .ZN(G1336gat));
  NOR2_X1   g587(.A1(new_n725), .A2(G92gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n778), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n783), .B2(new_n725), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n462), .A3(new_n786), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n794), .A2(G92gat), .B1(new_n778), .B2(new_n789), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n791), .ZN(G1337gat));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n575), .A3(new_n483), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n784), .A2(new_n736), .A3(new_n786), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n575), .ZN(G1338gat));
  OAI21_X1  g598(.A(G106gat), .B1(new_n783), .B2(new_n266), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n776), .A2(new_n777), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n266), .A2(G106gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n751), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n687), .A3(new_n786), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G106gat), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n804), .B(KEYINPUT109), .Z(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n776), .B2(new_n777), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n806), .B1(new_n813), .B2(KEYINPUT53), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n807), .B2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(KEYINPUT110), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n805), .B1(new_n814), .B2(new_n817), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n630), .A2(new_n632), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n633), .A2(KEYINPUT10), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n603), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n603), .B1(new_n633), .B2(KEYINPUT10), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n602), .B1(new_n820), .B2(new_n821), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n640), .B1(new_n828), .B2(new_n824), .ZN(new_n829));
  INV_X1    g628(.A(new_n635), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n827), .A2(new_n829), .B1(new_n830), .B2(new_n640), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n826), .B1(new_n634), .B2(new_n602), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n819), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n715), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n535), .B1(new_n534), .B2(new_n539), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n538), .A2(new_n545), .A3(new_n544), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n491), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n713), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n642), .A2(new_n643), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n693), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n598), .B2(new_n599), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n831), .A2(new_n834), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n707), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n658), .A2(new_n715), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n482), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n480), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n725), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n715), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n823), .A2(new_n627), .A3(new_n640), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n820), .A2(new_n825), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT55), .B1(new_n854), .B2(new_n828), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n822), .A2(new_n824), .A3(new_n603), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n641), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n852), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT55), .B1(new_n829), .B2(new_n832), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n693), .A3(new_n839), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n642), .A2(new_n643), .A3(new_n839), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n860), .B2(new_n715), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n693), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n846), .B1(new_n864), .B2(new_n707), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n462), .A2(new_n482), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR4_X1   g666(.A1(new_n865), .A2(new_n687), .A3(new_n443), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n554), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(G113gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n851), .B1(new_n868), .B2(new_n870), .ZN(G1340gat));
  INV_X1    g670(.A(G120gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n872), .A3(new_n751), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n868), .B2(new_n751), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(G1341gat));
  NAND2_X1  g678(.A1(new_n868), .A2(new_n657), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n707), .A2(G127gat), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n880), .A2(G127gat), .B1(new_n850), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT114), .Z(G1342gat));
  INV_X1    g682(.A(G134gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n868), .B2(new_n693), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT115), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n600), .A2(new_n462), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n848), .A2(new_n884), .A3(new_n849), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT56), .Z(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1343gat));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n266), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n858), .A2(new_n554), .A3(new_n859), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n600), .B1(new_n895), .B2(new_n862), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n844), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT117), .B(new_n600), .C1(new_n895), .C2(new_n862), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n657), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(new_n846), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT116), .B(new_n893), .C1(new_n865), .C2(new_n266), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n266), .B1(new_n845), .B2(new_n847), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(KEYINPUT57), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n736), .A2(new_n867), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n715), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G141gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n736), .A2(new_n266), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n554), .A2(G141gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n848), .A2(new_n725), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT118), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n892), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n892), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n906), .A2(new_n869), .A3(new_n907), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n891), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(G141gat), .ZN(new_n920));
  INV_X1    g719(.A(new_n916), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n913), .B1(new_n908), .B2(G141gat), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n922), .B(KEYINPUT119), .C1(new_n892), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n919), .A2(new_n924), .ZN(G1344gat));
  AND2_X1   g724(.A1(new_n848), .A2(new_n910), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n725), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n207), .A3(new_n751), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n906), .A2(new_n907), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n644), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(KEYINPUT59), .A3(new_n207), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n659), .A2(new_n554), .A3(new_n661), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n657), .B1(new_n896), .B2(new_n861), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT120), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n659), .A2(new_n554), .A3(new_n661), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n896), .A2(new_n861), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n657), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(new_n687), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n893), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n845), .A2(new_n847), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n894), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n751), .A3(new_n907), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n933), .B1(new_n946), .B2(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n929), .B1(new_n932), .B2(new_n947), .ZN(G1345gat));
  OAI21_X1  g747(.A(G155gat), .B1(new_n930), .B2(new_n707), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n928), .A2(new_n211), .A3(new_n657), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1346gat));
  OAI21_X1  g750(.A(G162gat), .B1(new_n930), .B2(new_n600), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n926), .A2(new_n212), .A3(new_n887), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n725), .A2(new_n664), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n849), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n715), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n955), .B(KEYINPUT121), .Z(new_n960));
  NOR4_X1   g759(.A1(new_n960), .A2(new_n865), .A3(new_n687), .A4(new_n443), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n554), .A2(new_n272), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1348gat));
  NAND3_X1  g762(.A1(new_n958), .A2(new_n273), .A3(new_n751), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n961), .A2(new_n751), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n273), .ZN(G1349gat));
  AOI21_X1  g765(.A(new_n310), .B1(new_n961), .B2(new_n657), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n957), .A2(new_n316), .A3(new_n707), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n969), .B(new_n970), .ZN(G1350gat));
  AOI21_X1  g770(.A(new_n291), .B1(new_n961), .B2(new_n693), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT61), .Z(new_n973));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n291), .A3(new_n693), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1351gat));
  AND2_X1   g774(.A1(new_n956), .A2(new_n910), .ZN(new_n976));
  AOI21_X1  g775(.A(G197gat), .B1(new_n976), .B2(new_n715), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n960), .A2(new_n736), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n942), .B2(new_n944), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n869), .A2(G197gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n982));
  XNOR2_X1  g781(.A(KEYINPUT123), .B(G204gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n976), .A2(new_n751), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n983), .B1(new_n979), .B2(new_n751), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n984), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n979), .A2(new_n751), .ZN(new_n990));
  INV_X1    g789(.A(new_n983), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n989), .A2(new_n992), .A3(KEYINPUT124), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n987), .A2(new_n993), .ZN(G1353gat));
  INV_X1    g793(.A(G211gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n995), .A3(new_n657), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n657), .ZN(new_n997));
  AND4_X1   g796(.A1(KEYINPUT125), .A2(new_n997), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n999));
  INV_X1    g798(.A(new_n999), .ZN(new_n1000));
  AOI22_X1  g799(.A1(new_n997), .A2(new_n1000), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n996), .B1(new_n998), .B2(new_n1001), .ZN(G1354gat));
  AOI21_X1  g801(.A(G218gat), .B1(new_n976), .B2(new_n693), .ZN(new_n1003));
  XOR2_X1   g802(.A(new_n1003), .B(KEYINPUT126), .Z(new_n1004));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005));
  OR2_X1    g804(.A1(new_n979), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n693), .A2(G218gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1007), .B1(new_n979), .B2(new_n1005), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1004), .B1(new_n1006), .B2(new_n1008), .ZN(G1355gat));
endmodule


