//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n210), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  AND3_X1   g0047(.A1(new_n247), .A2(KEYINPUT69), .A3(new_n213), .ZN(new_n248));
  AOI21_X1  g0048(.A(KEYINPUT69), .B1(new_n247), .B2(new_n213), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G13), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n214), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(G20), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G50), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(new_n250), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n214), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(G20), .B2(new_n203), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n256), .B1(G50), .B2(new_n257), .C1(new_n258), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n270), .A2(new_n272), .A3(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n272), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n273), .A2(G223), .B1(G77), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G222), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n275), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n290));
  AND2_X1   g0090(.A1(G1), .A2(G13), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT67), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(new_n251), .C1(G41), .C2(G45), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n289), .B1(new_n297), .B2(G226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n286), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n268), .B1(G190), .B2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n266), .A2(new_n267), .B1(new_n299), .B2(G200), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(new_n305), .A3(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n266), .B1(new_n300), .B2(G169), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n299), .A2(G179), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n281), .A2(new_n282), .A3(G232), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n282), .A2(G238), .A3(G1698), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n274), .A2(G107), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT70), .A4(new_n316), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n285), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n289), .B1(new_n297), .B2(G244), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n313), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n323), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(new_n324), .ZN(new_n331));
  INV_X1    g0131(.A(G77), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n259), .A2(new_n263), .B1(new_n214), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT15), .B(G87), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n260), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n250), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT72), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n254), .A2(G77), .A3(new_n255), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G77), .B2(new_n257), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n327), .A2(new_n331), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n312), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n259), .B1(new_n251), .B2(G20), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n254), .A2(new_n346), .B1(new_n253), .B2(new_n259), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT78), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n282), .B2(G20), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n271), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT7), .B(new_n214), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT77), .B1(new_n355), .B2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  INV_X1    g0157(.A(G68), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(new_n351), .C2(new_n354), .ZN(new_n359));
  INV_X1    g0159(.A(G58), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n358), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n361), .B2(new_n201), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n262), .A2(G159), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT16), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n356), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n358), .B1(new_n351), .B2(new_n354), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n250), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n349), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n274), .B2(new_n214), .ZN(new_n373));
  AOI211_X1 g0173(.A(new_n350), .B(G20), .C1(new_n270), .C2(new_n272), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n365), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n258), .B1(new_n376), .B2(new_n368), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n357), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n369), .A2(KEYINPUT77), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n364), .A2(new_n368), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(KEYINPUT78), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n348), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n282), .A2(G226), .A3(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  INV_X1    g0185(.A(G223), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n384), .B(new_n385), .C1(new_n283), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n285), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n289), .B1(new_n297), .B2(G232), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n330), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n389), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n313), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n345), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n367), .A2(new_n371), .A3(new_n349), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT78), .B1(new_n377), .B2(new_n381), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n347), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n394), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G190), .B2(new_n392), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n347), .C1(new_n396), .C2(new_n397), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n383), .A2(KEYINPUT17), .A3(new_n404), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n262), .A2(G50), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n411), .B(KEYINPUT76), .Z(new_n412));
  NOR2_X1   g0212(.A1(new_n260), .A2(new_n332), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(G20), .B2(new_n358), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n258), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n253), .A2(new_n358), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT12), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n254), .A2(G68), .A3(new_n255), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT68), .B(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(G226), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(new_n232), .B2(new_n277), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n282), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n293), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G238), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n296), .A2(new_n430), .B1(new_n432), .B2(new_n288), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n423), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n429), .B2(new_n433), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT75), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n281), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n428), .B1(new_n439), .B2(new_n274), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n285), .ZN(new_n441));
  INV_X1    g0241(.A(new_n433), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n435), .A3(new_n442), .ZN(new_n443));
  AND4_X1   g0243(.A1(KEYINPUT75), .A2(new_n437), .A3(new_n443), .A4(G190), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n422), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n435), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n429), .B2(new_n433), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n443), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT74), .B1(new_n448), .B2(G200), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT74), .ZN(new_n450));
  AOI211_X1 g0250(.A(new_n450), .B(new_n402), .C1(new_n447), .C2(new_n443), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n437), .A2(new_n443), .A3(G179), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n330), .B1(new_n447), .B2(new_n443), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT14), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n422), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(G190), .B1(new_n325), .B2(new_n326), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n329), .A2(G200), .A3(new_n324), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n340), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n344), .A2(new_n410), .A3(new_n461), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n251), .A2(G33), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n257), .B(new_n466), .C1(new_n248), .C2(new_n249), .ZN(new_n467));
  INV_X1    g0267(.A(G107), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n253), .A2(new_n468), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT25), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n270), .A2(new_n272), .A3(new_n214), .A4(G87), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT22), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n282), .A2(new_n476), .A3(new_n214), .A4(G87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n214), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n468), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT24), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n478), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n473), .B1(new_n490), .B2(new_n250), .ZN(new_n491));
  AOI211_X1 g0291(.A(KEYINPUT24), .B(new_n484), .C1(new_n475), .C2(new_n477), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n478), .B2(new_n485), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n473), .B(new_n250), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n472), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n270), .A2(new_n272), .A3(G257), .A4(G1698), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n282), .A2(KEYINPUT87), .A3(G257), .A4(G1698), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n281), .A2(new_n282), .A3(G250), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G294), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G41), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G1), .ZN(new_n508));
  INV_X1    g0308(.A(G41), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n293), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n503), .A2(new_n285), .B1(G264), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n431), .A2(new_n506), .A3(new_n508), .A4(new_n510), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n330), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n313), .A3(new_n515), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n496), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n472), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n250), .B1(new_n492), .B2(new_n493), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT86), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n524), .B2(new_n494), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n503), .A2(new_n285), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(G264), .ZN(new_n527));
  AND4_X1   g0327(.A1(G190), .A2(new_n526), .A3(new_n527), .A4(new_n515), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n402), .B1(new_n514), .B2(new_n515), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n282), .A2(G244), .A3(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n283), .C2(new_n430), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n285), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n293), .B(G250), .C1(G1), .C2(new_n507), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n431), .A2(new_n508), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n423), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n535), .B2(new_n285), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(G200), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n270), .A2(new_n272), .A3(new_n214), .A4(G68), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT83), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n282), .A2(new_n546), .A3(new_n214), .A4(G68), .ZN(new_n547));
  NOR3_X1   g0347(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n548));
  AOI21_X1  g0348(.A(G20), .B1(G33), .B2(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT19), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(new_n214), .A3(G33), .A4(G97), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n545), .A2(new_n547), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n553), .A2(KEYINPUT84), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(KEYINPUT84), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n250), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n253), .A2(new_n334), .ZN(new_n557));
  INV_X1    g0357(.A(new_n467), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G87), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n543), .A2(new_n556), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n542), .A2(G169), .ZN(new_n561));
  AOI211_X1 g0361(.A(G179), .B(new_n539), .C1(new_n535), .C2(new_n285), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n467), .A2(new_n334), .ZN(new_n564));
  INV_X1    g0364(.A(new_n555), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n250), .B1(new_n553), .B2(KEYINPUT84), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n557), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n355), .A2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n468), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT80), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT6), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n220), .A2(new_n468), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n572), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n262), .A2(G77), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT79), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n570), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n250), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT82), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n257), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n467), .B2(new_n220), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n582), .B1(new_n355), .B2(G107), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n258), .B1(new_n592), .B2(new_n580), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT82), .B1(new_n593), .B2(new_n589), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT4), .A4(G244), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G283), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  INV_X1    g0399(.A(G244), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n283), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n293), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n515), .B1(new_n512), .B2(new_n221), .ZN(new_n603));
  OAI21_X1  g0403(.A(G169), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n601), .A2(new_n596), .A3(new_n595), .A4(new_n597), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n285), .ZN(new_n606));
  INV_X1    g0406(.A(new_n603), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(G179), .A3(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n591), .A2(new_n594), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n585), .A2(new_n590), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n402), .B1(new_n606), .B2(new_n607), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n423), .B(new_n603), .C1(new_n605), .C2(new_n285), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n569), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT21), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n273), .A2(G264), .B1(G303), .B2(new_n274), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n281), .A2(new_n282), .A3(G257), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n293), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n511), .A2(G270), .A3(new_n293), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n515), .ZN(new_n620));
  OAI21_X1  g0420(.A(G169), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G116), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n467), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n247), .A2(new_n213), .B1(G20), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n596), .B(new_n214), .C1(G33), .C2(new_n220), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n624), .A2(KEYINPUT20), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT20), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(G20), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n626), .A2(new_n627), .B1(new_n252), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n615), .B1(new_n621), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n282), .A2(G264), .A3(G1698), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n274), .A2(G303), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n617), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n285), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n619), .A2(new_n515), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(G190), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n620), .B1(new_n285), .B2(new_n634), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n630), .B(new_n637), .C1(new_n402), .C2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n330), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(KEYINPUT21), .B1(new_n638), .B2(G179), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n631), .B(new_n639), .C1(new_n641), .C2(new_n630), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT85), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(G179), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n621), .B2(new_n615), .ZN(new_n646));
  INV_X1    g0446(.A(new_n630), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(KEYINPUT85), .A3(new_n631), .A4(new_n639), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n614), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n465), .A2(new_n532), .A3(new_n651), .ZN(G372));
  NAND2_X1  g0452(.A1(new_n407), .A2(new_n408), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(new_n453), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n460), .A2(new_n343), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n401), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n307), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n604), .A2(new_n608), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n586), .B1(new_n585), .B2(new_n590), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n593), .A2(KEYINPUT82), .A3(new_n589), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n569), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n557), .B(new_n559), .C1(new_n565), .C2(new_n566), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n664), .A2(new_n543), .B1(new_n567), .B2(new_n563), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n604), .A2(new_n608), .B1(new_n585), .B2(new_n590), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n662), .A2(new_n668), .A3(new_n568), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n648), .A2(new_n631), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT88), .B1(new_n496), .B2(new_n520), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n525), .A2(new_n672), .A3(new_n519), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n531), .A2(new_n665), .A3(new_n675), .A4(new_n661), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n669), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n311), .B(new_n657), .C1(new_n465), .C2(new_n678), .ZN(G369));
  OR3_X1    g0479(.A1(new_n252), .A2(KEYINPUT27), .A3(G20), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT27), .B1(new_n252), .B2(G20), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n644), .A2(new_n649), .B1(new_n647), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n684), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n670), .A2(new_n630), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT89), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n525), .A2(new_n686), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n532), .A2(KEYINPUT90), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT90), .B1(new_n532), .B2(new_n696), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n697), .B(new_n698), .C1(new_n521), .C2(new_n686), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n521), .A2(new_n672), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n524), .A2(new_n494), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n519), .B1(new_n702), .B2(new_n472), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT88), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n684), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n697), .A2(new_n698), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n670), .A2(new_n684), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n700), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n208), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n548), .A2(new_n622), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n211), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT93), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n678), .B2(new_n684), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n676), .B1(new_n705), .B2(new_n670), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT93), .B(new_n686), .C1(new_n720), .C2(new_n669), .ZN(new_n721));
  XOR2_X1   g0521(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n719), .A2(new_n721), .A3(KEYINPUT95), .A4(new_n722), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n676), .B1(new_n521), .B2(new_n670), .ZN(new_n728));
  INV_X1    g0528(.A(new_n667), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT26), .B1(new_n569), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n665), .A2(new_n666), .A3(new_n609), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n568), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n686), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n702), .A2(new_n530), .A3(new_n472), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n703), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n614), .A3(new_n650), .A4(new_n686), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT91), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n514), .A2(new_n740), .A3(new_n542), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n635), .A2(new_n636), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n313), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n740), .B1(new_n514), .B2(new_n542), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n603), .B1(new_n605), .B2(new_n285), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT30), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n514), .A2(new_n542), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n602), .A2(new_n751), .A3(new_n603), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n750), .A2(new_n752), .A3(new_n743), .A4(new_n741), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n638), .A2(new_n542), .A3(G179), .ZN(new_n754));
  INV_X1    g0554(.A(new_n747), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n754), .A2(new_n516), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n684), .B1(new_n748), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n744), .A2(new_n755), .A3(new_n745), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n753), .B(new_n756), .C1(new_n761), .C2(KEYINPUT30), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n739), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n764), .A2(KEYINPUT92), .A3(G330), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT92), .B1(new_n764), .B2(G330), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n736), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n717), .B1(new_n768), .B2(G1), .ZN(G364));
  INV_X1    g0569(.A(new_n695), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n214), .A2(G13), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n771), .A2(KEYINPUT96), .A3(new_n507), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n251), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT96), .B1(new_n771), .B2(new_n507), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n712), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n688), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n770), .B(new_n777), .C1(G330), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n214), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  AOI21_X1  g0582(.A(new_n213), .B1(G20), .B2(new_n330), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT98), .Z(new_n786));
  NAND3_X1  g0586(.A1(new_n208), .A2(G355), .A3(new_n282), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G116), .B2(new_n208), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n242), .A2(new_n507), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n208), .A2(new_n274), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n507), .B2(new_n212), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n776), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n423), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n313), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n220), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n214), .A2(new_n313), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n423), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n202), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(G190), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n798), .B(new_n803), .C1(G68), .C2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n799), .A2(new_n423), .A3(new_n402), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n282), .B1(new_n806), .B2(new_n332), .ZN(new_n807));
  NOR4_X1   g0607(.A1(new_n214), .A2(new_n423), .A3(new_n402), .A4(G179), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(G87), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n423), .A2(G20), .ZN(new_n810));
  AOI21_X1  g0610(.A(G179), .B1(new_n810), .B2(KEYINPUT100), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(KEYINPUT100), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n402), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G107), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n799), .A2(new_n794), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G58), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n805), .A2(new_n809), .A3(new_n814), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n812), .A2(G200), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G159), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n826));
  XNOR2_X1  g0626(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n274), .B1(new_n806), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G303), .B2(new_n808), .ZN(new_n830));
  INV_X1    g0630(.A(new_n804), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT33), .B(G317), .Z(new_n832));
  INV_X1    g0632(.A(G322), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n833), .C2(new_n820), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n801), .A2(G326), .B1(new_n796), .B2(G294), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(KEYINPUT102), .B1(new_n813), .B2(G283), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n824), .A2(G329), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(KEYINPUT102), .C2(new_n835), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n823), .A2(new_n827), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n793), .B1(new_n839), .B2(new_n783), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n778), .B2(new_n782), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n779), .A2(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n341), .A2(new_n684), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n464), .A2(new_n342), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT107), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n343), .A2(new_n684), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT107), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n464), .A2(new_n342), .A3(new_n847), .A4(new_n843), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n719), .A2(new_n721), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n674), .A2(new_n677), .ZN(new_n852));
  INV_X1    g0652(.A(new_n669), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n684), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n845), .A2(new_n848), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n776), .B1(new_n857), .B2(new_n767), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n767), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n783), .A2(new_n780), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n808), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n274), .B1(new_n862), .B2(new_n468), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n798), .B(new_n863), .C1(new_n821), .C2(G294), .ZN(new_n864));
  INV_X1    g0664(.A(new_n824), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n828), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n806), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G303), .A2(new_n801), .B1(new_n867), .B2(G116), .ZN(new_n868));
  INV_X1    g0668(.A(G283), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n831), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT103), .Z(new_n871));
  AOI211_X1 g0671(.A(new_n866), .B(new_n871), .C1(G87), .C2(new_n813), .ZN(new_n872));
  AOI22_X1  g0672(.A1(G137), .A2(new_n801), .B1(new_n804), .B2(G150), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT104), .Z(new_n874));
  INV_X1    g0674(.A(G143), .ZN(new_n875));
  INV_X1    g0675(.A(G159), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n874), .B1(new_n875), .B2(new_n820), .C1(new_n876), .C2(new_n806), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT34), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n274), .B1(new_n824), .B2(G132), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT105), .Z(new_n880));
  NAND2_X1  g0680(.A1(new_n813), .A2(G68), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n881), .B1(new_n202), .B2(new_n862), .C1(new_n360), .C2(new_n797), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n872), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n776), .B1(G77), .B2(new_n861), .C1(new_n884), .C2(new_n784), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT106), .Z(new_n886));
  INV_X1    g0686(.A(new_n780), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n849), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n859), .A2(new_n888), .ZN(G384));
  OR2_X1    g0689(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(G116), .A3(new_n215), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT36), .Z(new_n893));
  OR3_X1    g0693(.A1(new_n361), .A2(new_n211), .A3(new_n332), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n202), .A2(G68), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n251), .B(G13), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n739), .A2(new_n763), .ZN(new_n898));
  AOI211_X1 g0698(.A(KEYINPUT111), .B(KEYINPUT31), .C1(new_n762), .C2(new_n684), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT111), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n758), .B2(new_n759), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n465), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n739), .B(new_n763), .C1(new_n899), .C2(new_n901), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n422), .A2(new_n686), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n453), .B2(new_n460), .ZN(new_n907));
  INV_X1    g0707(.A(new_n459), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n421), .B1(new_n908), .B2(new_n457), .ZN(new_n909));
  INV_X1    g0709(.A(new_n906), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(new_n452), .C2(new_n445), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(new_n849), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n392), .A2(G169), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(new_n682), .C1(new_n313), .C2(new_n392), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n398), .A2(new_n917), .ZN(new_n918));
  AND4_X1   g0718(.A1(KEYINPUT110), .A2(new_n918), .A3(KEYINPUT37), .A4(new_n405), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT110), .ZN(new_n920));
  INV_X1    g0720(.A(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n383), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .B1(new_n918), .B2(new_n405), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n383), .A2(new_n682), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n395), .A2(new_n400), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n653), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n915), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n356), .A2(new_n359), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT16), .B1(new_n929), .B2(new_n365), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n381), .A2(new_n250), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n347), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n682), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n407), .A2(new_n408), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n401), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n917), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n405), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT37), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT37), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n918), .A2(new_n940), .A3(new_n405), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT38), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n936), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n905), .B(new_n913), .C1(new_n928), .C2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n936), .B2(new_n942), .ZN(new_n946));
  INV_X1    g0746(.A(new_n934), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n926), .B2(new_n653), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n939), .A2(new_n941), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(KEYINPUT38), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT40), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n912), .A2(new_n849), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n902), .B2(new_n898), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n945), .A2(KEYINPUT40), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n904), .B1(new_n954), .B2(new_n689), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n924), .A2(new_n927), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n409), .A2(new_n947), .B1(new_n939), .B2(new_n941), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n959), .A2(new_n914), .B1(new_n960), .B2(KEYINPUT38), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n913), .A2(new_n905), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT40), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n951), .A2(new_n953), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n957), .B(new_n958), .C1(new_n965), .C2(new_n903), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n460), .A2(new_n686), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT108), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT38), .B1(new_n948), .B2(new_n949), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(KEYINPUT39), .C1(new_n944), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n959), .A2(new_n914), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT39), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n950), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n946), .A2(new_n950), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n969), .B1(new_n976), .B2(KEYINPUT39), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n968), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n342), .A2(new_n684), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n854), .B2(new_n855), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n976), .A3(new_n912), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n926), .A2(new_n682), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n657), .A2(new_n311), .ZN(new_n986));
  INV_X1    g0786(.A(new_n735), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n465), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n727), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n985), .B(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n966), .A2(new_n990), .B1(G1), .B2(new_n771), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT113), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n991), .A2(new_n992), .B1(new_n990), .B2(new_n966), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n897), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT114), .Z(G367));
  INV_X1    g0796(.A(new_n238), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n997), .A2(new_n790), .B1(new_n208), .B2(new_n334), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n797), .A2(new_n358), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n831), .A2(new_n876), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G143), .C2(new_n801), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n282), .B1(new_n202), .B2(new_n806), .C1(new_n862), .C2(new_n360), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n821), .B2(G150), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n824), .A2(G137), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n813), .A2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n808), .A2(G116), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT46), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n274), .B1(new_n869), .B2(new_n806), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G303), .B2(new_n821), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1007), .A2(new_n1008), .B1(new_n801), .B2(G311), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n804), .A2(G294), .B1(new_n796), .B2(G107), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n813), .A2(G97), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n865), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1006), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n776), .B1(new_n786), .B2(new_n998), .C1(new_n1018), .C2(new_n784), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT118), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n663), .A2(new_n684), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT115), .Z(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n567), .A3(new_n563), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n569), .B2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1020), .B1(new_n782), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT116), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n707), .A2(new_n708), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n610), .A2(new_n684), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n675), .A2(new_n661), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n667), .A2(new_n684), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT42), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT42), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n661), .B1(new_n1033), .B2(new_n521), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n686), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1034), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT43), .B2(new_n1024), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1040), .A2(KEYINPUT43), .A3(new_n1024), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n700), .A2(new_n1033), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1027), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1043), .A2(KEYINPUT116), .A3(new_n1046), .A4(new_n1044), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n775), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n768), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n709), .A2(new_n1032), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT45), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT45), .B1(new_n709), .B2(new_n1032), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OR3_X1    g0858(.A1(new_n709), .A2(KEYINPUT44), .A3(new_n1032), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT44), .B1(new_n709), .B2(new_n1032), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT117), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n700), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n700), .A2(new_n1063), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n695), .A2(KEYINPUT117), .A3(new_n699), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1065), .A2(new_n1058), .A3(new_n1066), .A4(new_n1061), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1028), .B1(new_n699), .B2(new_n708), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n695), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1053), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n712), .B(KEYINPUT41), .Z(new_n1072));
  OAI21_X1  g0872(.A(new_n1052), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1026), .B1(new_n1051), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G387));
  OR2_X1    g0875(.A1(new_n768), .A2(new_n1070), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n768), .A2(new_n1070), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n712), .B(KEYINPUT121), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n699), .A2(new_n782), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n786), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n468), .B2(new_n208), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n235), .A2(G45), .A3(new_n274), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT50), .B1(new_n259), .B2(G50), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n507), .C1(new_n358), .C2(new_n332), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n259), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n274), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n714), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n711), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n776), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n797), .A2(new_n334), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n259), .B2(new_n831), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G159), .B2(new_n801), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n282), .B1(new_n358), .B2(new_n806), .C1(new_n862), .C2(new_n332), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n821), .B2(G50), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n824), .A2(G150), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1014), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G294), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n797), .A2(new_n869), .B1(new_n862), .B2(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n831), .A2(new_n828), .B1(new_n802), .B2(new_n833), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT120), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(KEYINPUT120), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n821), .A2(G317), .B1(G303), .B2(new_n867), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT48), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1100), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT49), .Z(new_n1109));
  AOI21_X1  g0909(.A(new_n282), .B1(new_n824), .B2(G326), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n813), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n622), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1098), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1090), .B1(new_n1113), .B2(new_n783), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1070), .A2(new_n775), .B1(new_n1080), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1079), .A2(new_n1115), .ZN(G393));
  INV_X1    g0916(.A(new_n1078), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1077), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n1068), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1118), .B2(new_n1068), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1068), .A2(new_n775), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1032), .A2(new_n782), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n790), .A2(new_n245), .B1(new_n220), .B2(new_n208), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n776), .B1(new_n786), .B2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n831), .A2(new_n202), .B1(new_n797), .B2(new_n332), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n282), .B1(new_n259), .B2(new_n806), .C1(new_n862), .C2(new_n358), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(G87), .C2(new_n813), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n875), .B2(new_n865), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n820), .A2(new_n876), .B1(new_n261), .B2(new_n802), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT51), .Z(new_n1130));
  OAI22_X1  g0930(.A1(new_n820), .A2(new_n828), .B1(new_n1015), .B2(new_n802), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT52), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n824), .A2(G322), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n274), .B1(new_n806), .B2(new_n1099), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G283), .B2(new_n808), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n804), .A2(G303), .B1(new_n796), .B2(G116), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n814), .A2(new_n1133), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1128), .A2(new_n1130), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1124), .B1(new_n1138), .B2(new_n783), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1122), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1121), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1120), .A2(new_n1141), .ZN(G390));
  AND2_X1   g0942(.A1(new_n849), .A2(G330), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1143), .A2(new_n905), .A3(new_n912), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT39), .B1(new_n944), .B2(new_n970), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT108), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n912), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n967), .B1(new_n980), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1147), .A2(new_n974), .A3(new_n971), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n855), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n733), .A2(new_n1151), .B1(new_n342), .B2(new_n684), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n912), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n967), .C1(new_n944), .C2(new_n928), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1145), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n849), .B(new_n912), .C1(new_n765), .C2(new_n766), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1143), .A2(new_n905), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1152), .B1(new_n1160), .B2(new_n1148), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1157), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n849), .B1(new_n765), .B2(new_n766), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1144), .B1(new_n1163), .B2(new_n1148), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n980), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n989), .A3(new_n904), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1159), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n989), .A2(new_n904), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1169), .A2(new_n1156), .A3(new_n1158), .A4(new_n1165), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1170), .A3(new_n1078), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT54), .B(G143), .Z(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT122), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n867), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G128), .A2(new_n801), .B1(new_n804), .B2(G137), .ZN(new_n1175));
  INV_X1    g0975(.A(G132), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1174), .B(new_n1175), .C1(new_n1176), .C2(new_n820), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n824), .A2(G125), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n862), .A2(KEYINPUT53), .A3(new_n261), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT53), .B1(new_n862), .B2(new_n261), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n876), .B2(new_n797), .ZN(new_n1181));
  OR4_X1    g0981(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n274), .B1(new_n813), .B2(G50), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(KEYINPUT123), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(KEYINPUT123), .B2(new_n1183), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n797), .A2(new_n332), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n802), .A2(new_n869), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G107), .C2(new_n804), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n274), .B1(new_n220), .B2(new_n806), .C1(new_n862), .C2(new_n218), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n821), .B2(G116), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n824), .A2(G294), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1190), .A3(new_n881), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n784), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n777), .B(new_n1193), .C1(new_n259), .C2(new_n860), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT124), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1147), .A2(new_n974), .A3(new_n971), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1197), .B2(new_n780), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1159), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n775), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1171), .A2(new_n1200), .ZN(G378));
  AND3_X1   g1001(.A1(new_n1150), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1166), .A2(new_n1202), .A3(new_n1155), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1168), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n982), .A2(new_n983), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1196), .B2(new_n968), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1207));
  NAND2_X1  g1007(.A1(new_n312), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n266), .A2(new_n933), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT125), .Z(new_n1210));
  AOI21_X1  g1010(.A(new_n310), .B1(new_n304), .B2(new_n306), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1207), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1210), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n310), .B(new_n1207), .C1(new_n304), .C2(new_n306), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n965), .B2(G330), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n689), .B(new_n1219), .C1(new_n963), .C2(new_n964), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1206), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1219), .B1(new_n954), .B2(new_n689), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n965), .A2(G330), .A3(new_n1220), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n985), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT126), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1206), .B(KEYINPUT126), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1078), .B1(new_n1204), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1170), .A2(new_n1169), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1219), .A2(new_n887), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n821), .A2(G128), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G137), .A2(new_n867), .B1(new_n796), .B2(G150), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G125), .A2(new_n801), .B1(new_n804), .B2(G132), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1173), .A2(new_n808), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n269), .B(new_n509), .C1(new_n1111), .C2(new_n876), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G124), .B2(new_n824), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1111), .A2(new_n360), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n831), .A2(new_n220), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n999), .B(new_n1248), .C1(G116), .C2(new_n801), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n282), .A2(G41), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n334), .B2(new_n806), .C1(new_n862), .C2(new_n332), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n821), .B2(G107), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1247), .B(new_n1253), .C1(G283), .C2(new_n824), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1250), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1257), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1258));
  AND4_X1   g1058(.A1(new_n1246), .A2(new_n1255), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n776), .B1(G50), .B2(new_n861), .C1(new_n1259), .C2(new_n784), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1236), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1233), .B2(new_n775), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1235), .A2(new_n1262), .ZN(G375));
  INV_X1    g1063(.A(new_n1165), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1168), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1072), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1166), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n274), .B1(new_n468), .B2(new_n806), .C1(new_n862), .C2(new_n220), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1092), .B1(new_n831), .B2(new_n622), .C1(new_n1099), .C2(new_n802), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(G283), .C2(new_n821), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G77), .A2(new_n813), .B1(new_n824), .B2(G303), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n821), .A2(G137), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n282), .B1(new_n261), .B2(new_n806), .C1(new_n862), .C2(new_n876), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1173), .A2(new_n804), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n802), .A2(new_n1176), .B1(new_n797), .B2(new_n202), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1247), .B1(G128), .B2(new_n824), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1270), .A2(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n776), .B1(G68), .B2(new_n861), .C1(new_n1278), .C2(new_n784), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1148), .B2(new_n780), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1165), .B2(new_n775), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1267), .A2(new_n1281), .ZN(G381));
  NOR2_X1   g1082(.A1(G390), .A2(G384), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1171), .A2(new_n1200), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1079), .A2(new_n779), .A3(new_n841), .A4(new_n1115), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1285), .A2(G381), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1287), .A2(G375), .A3(G387), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1288), .B(new_n1289), .ZN(G407));
  NOR3_X1   g1090(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1291));
  INV_X1    g1091(.A(G213), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G407), .A2(new_n1293), .ZN(G409));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1262), .C1(new_n1231), .C2(new_n1234), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1266), .B(new_n1233), .C1(new_n1203), .C2(new_n1168), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1261), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1297), .B(new_n1298), .C1(new_n1052), .C2(new_n1230), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1284), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1292), .A2(G343), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT60), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1265), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1168), .A2(new_n1264), .A3(KEYINPUT60), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1306), .A2(new_n1078), .A3(new_n1166), .A4(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1308), .A2(G384), .A3(new_n1281), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G384), .B1(new_n1308), .B2(new_n1281), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1295), .B1(new_n1304), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G393), .A2(G396), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1285), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n1120), .A3(new_n1141), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(G390), .A2(new_n1285), .A3(new_n1314), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1316), .A2(new_n1074), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1074), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G2897), .B(new_n1302), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1310), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1308), .A2(G384), .A3(new_n1281), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1302), .A2(G2897), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1304), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1302), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1311), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1313), .A2(new_n1320), .A3(new_n1327), .A4(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1328), .A2(new_n1331), .A3(new_n1311), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1333), .B1(new_n1328), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1331), .B1(new_n1328), .B2(new_n1311), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1332), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1330), .B1(new_n1337), .B2(new_n1320), .ZN(G405));
  AOI21_X1  g1138(.A(G378), .B1(new_n1235), .B2(new_n1262), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1296), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1311), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1339), .A2(new_n1311), .A3(new_n1340), .ZN(new_n1343));
  OAI22_X1  g1143(.A1(new_n1342), .A2(new_n1343), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1343), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(new_n1320), .A3(new_n1341), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(G402));
endmodule


