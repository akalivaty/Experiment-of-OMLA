//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G244), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n218), .A2(G77), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(new_n206), .A2(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G50), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  INV_X1    g0047(.A(G13), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n248), .A2(new_n207), .A3(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n248), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n247), .A2(new_n253), .B1(G50), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n251), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT8), .B(G58), .Z(new_n258));
  NAND2_X1  g0058(.A1(new_n207), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(new_n260), .B1(G150), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n203), .A2(G20), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT9), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G274), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n273), .B1(G226), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G222), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(new_n274), .C1(G77), .C2(new_n281), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n277), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(G200), .A3(new_n290), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n267), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n267), .A2(new_n292), .A3(new_n298), .A4(new_n293), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n296), .A2(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n229), .A2(G1698), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n281), .B(new_n303), .C1(G226), .C2(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n270), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(G238), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n274), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n275), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n317), .A3(G169), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n313), .B1(new_n306), .B2(new_n311), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n320), .C1(KEYINPUT73), .C2(new_n312), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G68), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n249), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n259), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n252), .A2(G68), .A3(new_n245), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT11), .B1(new_n329), .B2(new_n251), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n323), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n314), .B2(G200), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n321), .A2(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n291), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n265), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n289), .A2(new_n343), .A3(new_n290), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n273), .B1(new_n218), .B2(new_n276), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n347), .B(KEYINPUT69), .Z(new_n348));
  NAND3_X1  g0148(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n281), .A2(G232), .A3(new_n283), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT70), .B(G107), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n350), .C1(new_n281), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n274), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n252), .A2(G77), .A3(new_n245), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G77), .B2(new_n255), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n258), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n259), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n251), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n355), .B(new_n361), .C1(new_n362), .C2(new_n354), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n361), .B1(new_n354), .B2(new_n343), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n348), .A2(new_n340), .A3(new_n353), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n302), .A2(new_n339), .A3(new_n346), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n258), .A2(new_n245), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n253), .A2(new_n369), .B1(new_n255), .B2(new_n258), .ZN(new_n370));
  INV_X1    g0170(.A(G58), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n324), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n201), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n261), .A2(G159), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(KEYINPUT16), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AND2_X1   g0177(.A1(KEYINPUT74), .A2(G33), .ZN(new_n378));
  NOR2_X1   g0178(.A1(KEYINPUT74), .A2(G33), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n378), .A2(new_n379), .A3(new_n278), .ZN(new_n380));
  INV_X1    g0180(.A(new_n279), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n377), .B(new_n207), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G68), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT74), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n268), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT74), .A2(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT3), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n279), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n377), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n376), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT75), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n324), .B1(new_n388), .B2(new_n377), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n378), .A2(new_n379), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n381), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT7), .B1(new_n394), .B2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT75), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n376), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n257), .B1(new_n391), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n377), .A2(G20), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT77), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n280), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT74), .B(G33), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n403), .A3(new_n278), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n401), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n279), .A2(new_n280), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(new_n207), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n324), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n373), .A2(new_n374), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n400), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n370), .B1(new_n399), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n270), .A2(G232), .A3(new_n272), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n310), .ZN(new_n418));
  MUX2_X1   g0218(.A(G223), .B(G226), .S(G1698), .Z(new_n419));
  NAND2_X1  g0219(.A1(new_n394), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n270), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n418), .A2(new_n340), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n422), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n416), .A2(KEYINPUT78), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(KEYINPUT78), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n273), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n343), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT18), .B1(new_n415), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n370), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n397), .B1(new_n396), .B2(new_n376), .ZN(new_n432));
  AOI211_X1 g0232(.A(KEYINPUT75), .B(new_n375), .C1(new_n392), .C2(new_n395), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n251), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n400), .ZN(new_n435));
  INV_X1    g0235(.A(new_n401), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n405), .A2(new_n278), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(KEYINPUT77), .B1(KEYINPUT3), .B2(new_n268), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n438), .B2(new_n406), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n439), .B2(new_n410), .ZN(new_n440));
  INV_X1    g0240(.A(new_n413), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n431), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  INV_X1    g0244(.A(new_n429), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n430), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G200), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n418), .B2(new_n422), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n424), .A2(new_n427), .A3(new_n362), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n431), .B(new_n451), .C1(new_n434), .C2(new_n442), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n399), .A2(new_n414), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n431), .A4(new_n451), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n368), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n387), .A2(new_n279), .ZN(new_n463));
  INV_X1    g0263(.A(G257), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n463), .A2(new_n464), .A3(new_n283), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT89), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n394), .A2(G257), .A3(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT89), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n394), .A2(G250), .A3(new_n283), .ZN(new_n471));
  XOR2_X1   g0271(.A(KEYINPUT90), .B(G294), .Z(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n405), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n274), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT5), .B(G41), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n271), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n270), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n477), .A2(G190), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n474), .B1(new_n467), .B2(new_n469), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n483), .B(new_n486), .C1(new_n488), .C2(new_n270), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT87), .B1(new_n255), .B2(G107), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n249), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(KEYINPUT25), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n252), .B1(G1), .B2(new_n268), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT25), .B1(new_n491), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT88), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n251), .B(new_n249), .C1(new_n206), .C2(G33), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(new_n498), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT88), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n495), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n394), .A2(KEYINPUT22), .A3(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n405), .A2(G116), .ZN(new_n507));
  AOI21_X1  g0307(.A(G20), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n351), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT23), .B1(new_n509), .B2(new_n207), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n409), .A2(G20), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n510), .B(new_n511), .C1(new_n513), .C2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n508), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n508), .B2(new_n514), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n251), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n487), .A2(new_n490), .A3(new_n505), .A4(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n477), .A2(new_n340), .A3(new_n483), .A4(new_n486), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n489), .A2(new_n343), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n251), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n505), .B1(new_n523), .B2(new_n516), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT91), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n520), .A2(new_n525), .A3(KEYINPUT91), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n394), .A2(new_n207), .A3(G68), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  INV_X1    g0332(.A(G97), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n351), .A2(new_n512), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n305), .A2(new_n207), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n259), .A2(KEYINPUT19), .A3(new_n533), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n251), .B1(new_n249), .B2(new_n359), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n500), .A2(G87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n309), .A2(new_n480), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n270), .B(G250), .C1(G1), .C2(new_n479), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  MUX2_X1   g0348(.A(G238), .B(G244), .S(G1698), .Z(new_n549));
  NAND2_X1  g0349(.A1(new_n394), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n270), .B1(new_n550), .B2(new_n507), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n448), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT84), .B1(new_n541), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n543), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT82), .B1(new_n542), .B2(new_n543), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(G200), .B1(new_n557), .B2(new_n551), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT84), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n539), .A4(new_n540), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n557), .A2(new_n551), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G190), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n554), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n561), .A2(new_n343), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n548), .A2(new_n552), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n340), .ZN(new_n566));
  INV_X1    g0366(.A(new_n359), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n500), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n539), .A2(KEYINPUT83), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT83), .B1(new_n539), .B2(new_n568), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n564), .A2(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT85), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n563), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n563), .B2(new_n571), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  INV_X1    g0375(.A(G270), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n483), .B1(new_n576), .B2(new_n484), .ZN(new_n577));
  MUX2_X1   g0377(.A(G257), .B(G264), .S(G1698), .Z(new_n578));
  AOI22_X1  g0378(.A1(new_n394), .A2(new_n578), .B1(G303), .B2(new_n409), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n270), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G283), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n582), .B(new_n207), .C1(G33), .C2(new_n533), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(new_n251), .C1(new_n207), .C2(G116), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n584), .B(KEYINPUT20), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT86), .B1(new_n255), .B2(G116), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n249), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n496), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(G169), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n575), .B1(new_n581), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(G200), .B1(new_n577), .B2(new_n580), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n482), .B1(new_n485), .B2(G270), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(G190), .C1(new_n270), .C2(new_n579), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n585), .A2(new_n591), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n591), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n584), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n595), .B1(new_n270), .B2(new_n579), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT21), .A4(G169), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n581), .A2(new_n602), .A3(G179), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n593), .A2(new_n598), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n351), .B1(new_n408), .B2(new_n411), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n261), .A2(G77), .ZN(new_n608));
  XNOR2_X1  g0408(.A(G97), .B(G107), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT80), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(KEYINPUT6), .ZN(new_n611));
  MUX2_X1   g0411(.A(new_n610), .B(G97), .S(KEYINPUT6), .Z(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n608), .B1(new_n613), .B2(new_n207), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n251), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n255), .A2(G97), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n500), .B2(G97), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n619), .A2(new_n620), .A3(new_n582), .ZN(new_n621));
  XOR2_X1   g0421(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n622));
  NAND2_X1  g0422(.A1(new_n283), .A2(G244), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n463), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n270), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n483), .B1(new_n464), .B2(new_n484), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n340), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n343), .B1(new_n625), .B2(new_n626), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n618), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(G190), .ZN(new_n631));
  OAI21_X1  g0431(.A(G200), .B1(new_n625), .B2(new_n626), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n631), .A2(new_n615), .A3(new_n617), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n606), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n573), .A2(new_n574), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n462), .A2(new_n530), .A3(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n574), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n563), .A2(new_n571), .A3(new_n572), .ZN(new_n638));
  INV_X1    g0438(.A(new_n630), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n539), .A2(new_n568), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n564), .B2(new_n566), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT92), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n562), .A2(new_n539), .A3(new_n558), .A4(new_n540), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n639), .A2(new_n644), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n593), .A2(new_n604), .A3(new_n605), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n522), .A2(new_n524), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n520), .A2(new_n650), .B1(new_n651), .B2(new_n521), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n630), .A2(new_n644), .A3(new_n633), .A4(new_n648), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n646), .B(new_n649), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n462), .B1(new_n642), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n415), .A2(KEYINPUT18), .A3(new_n429), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n338), .A2(new_n365), .A3(new_n364), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n335), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n457), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n296), .A2(new_n297), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n300), .A2(new_n301), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n346), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n655), .A2(new_n665), .ZN(G369));
  NAND2_X1  g0466(.A1(new_n254), .A2(new_n207), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(G213), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n597), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT94), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n606), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n675), .B2(new_n606), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n650), .A2(new_n674), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n525), .A2(new_n673), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n524), .A2(new_n672), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n530), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n530), .A2(new_n650), .A3(new_n673), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n651), .A2(new_n521), .A3(new_n673), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n210), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n534), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n213), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  INV_X1    g0497(.A(new_n654), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n672), .B1(new_n698), .B2(new_n641), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n644), .A2(new_n648), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT26), .B1(new_n702), .B2(new_n630), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n703), .B(new_n646), .C1(new_n652), .C2(new_n653), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n637), .A2(new_n647), .A3(new_n638), .A4(new_n639), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n672), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n635), .A2(new_n530), .A3(new_n673), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n477), .A2(new_n486), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n603), .A2(new_n340), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n565), .A2(new_n625), .A3(new_n626), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(KEYINPUT30), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n627), .A2(G179), .A3(new_n581), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT95), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n565), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n561), .A2(KEYINPUT95), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n717), .A2(new_n489), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n627), .A3(new_n561), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n477), .A2(new_n486), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n716), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n726), .B2(new_n672), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n711), .B1(new_n712), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n710), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n697), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n681), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n248), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n206), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n692), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G330), .B2(new_n680), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n215), .B1(G20), .B2(new_n343), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n207), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(G303), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(new_n340), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n749), .A2(new_n362), .A3(new_n448), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G326), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n409), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n362), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n207), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n747), .B(new_n753), .C1(new_n472), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n744), .A2(new_n362), .A3(G200), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G283), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n749), .A2(new_n448), .A3(G190), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n749), .A2(new_n362), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G322), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n748), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n770), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n744), .A2(new_n772), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G329), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n757), .A2(new_n763), .A3(new_n768), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n764), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n780), .A2(new_n324), .B1(new_n751), .B2(new_n202), .ZN(new_n781));
  INV_X1    g0581(.A(new_n773), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G77), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n762), .A2(G107), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n755), .A2(new_n533), .ZN(new_n787));
  INV_X1    g0587(.A(new_n745), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n786), .B(new_n787), .C1(G87), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT32), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n777), .B2(G159), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n409), .B(new_n791), .C1(G58), .C2(new_n769), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n783), .A2(new_n784), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n743), .B1(new_n779), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n248), .A2(new_n268), .A3(KEYINPUT97), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT97), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G13), .B2(G33), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n742), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n210), .A2(new_n281), .ZN(new_n803));
  INV_X1    g0603(.A(G355), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(G116), .B2(new_n210), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n243), .A2(G45), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n691), .A2(new_n394), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(G45), .C2(new_n213), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n802), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n739), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n794), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n800), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n680), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n741), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  AOI22_X1  g0616(.A1(new_n764), .A2(G150), .B1(G159), .B2(new_n782), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n751), .C1(new_n819), .C2(new_n770), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT34), .Z(new_n821));
  AOI22_X1  g0621(.A1(new_n756), .A2(G58), .B1(new_n788), .B2(G50), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n463), .B1(G132), .B2(new_n777), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(new_n761), .C2(new_n324), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n780), .A2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n751), .A2(new_n746), .B1(new_n776), .B2(new_n774), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G294), .C2(new_n769), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n281), .B(new_n787), .C1(G116), .C2(new_n782), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n493), .C2(new_n745), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n761), .A2(new_n512), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n821), .A2(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n742), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n798), .A2(new_n742), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n739), .C1(G77), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n363), .B1(new_n361), .B2(new_n673), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n366), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n366), .A2(new_n672), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n836), .B1(new_n841), .B2(new_n798), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n700), .A2(new_n841), .ZN(new_n843));
  INV_X1    g0643(.A(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n699), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n739), .B1(new_n846), .B2(new_n731), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(new_n730), .A3(new_n845), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  OAI21_X1  g0650(.A(new_n462), .B1(new_n701), .B2(new_n709), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n665), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT104), .Z(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n415), .B2(new_n670), .ZN(new_n856));
  INV_X1    g0656(.A(new_n670), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n443), .A2(KEYINPUT101), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n452), .B(new_n860), .C1(new_n415), .C2(new_n429), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n391), .A2(new_n398), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n396), .A2(new_n441), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n257), .B1(new_n865), .B2(new_n400), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n370), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n863), .B1(new_n867), .B2(new_n670), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n432), .A2(new_n433), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n413), .B1(new_n392), .B2(new_n395), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n251), .B1(new_n870), .B2(new_n435), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n431), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(KEYINPUT100), .A3(new_n857), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n445), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n868), .A2(new_n873), .A3(new_n452), .A4(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n859), .A2(new_n862), .B1(new_n875), .B2(KEYINPUT37), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n868), .A2(new_n873), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n454), .A2(new_n456), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n658), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n854), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n868), .A2(new_n873), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n447), .B2(new_n457), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n861), .B1(new_n856), .B2(new_n858), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT38), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT102), .B(new_n854), .C1(new_n876), .C2(new_n879), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n443), .A2(new_n445), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n452), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n860), .B1(new_n893), .B2(new_n859), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n458), .B2(new_n859), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n885), .A2(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT39), .B1(new_n897), .B2(new_n886), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n890), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n335), .A2(new_n672), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n887), .B2(new_n888), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT103), .B1(new_n903), .B2(new_n898), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n845), .A2(new_n840), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n339), .A2(new_n334), .A3(new_n672), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n334), .A2(new_n672), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n335), .A2(new_n338), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n905), .B1(new_n658), .B2(new_n857), .C1(new_n889), .C2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n853), .B(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n897), .ZN(new_n914));
  INV_X1    g0714(.A(new_n886), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n712), .A2(new_n729), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n844), .A3(new_n910), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT40), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n918), .A2(KEYINPUT40), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n920), .B2(new_n889), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n462), .A2(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n921), .A2(new_n922), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n925), .A3(new_n711), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n913), .A2(new_n926), .B1(new_n206), .B2(new_n736), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n913), .B2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  OAI211_X1 g0729(.A(G116), .B(new_n216), .C1(new_n613), .C2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n613), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n214), .B(G77), .C1(new_n371), .C2(new_n324), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n202), .A2(G68), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n206), .B(G13), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n928), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n639), .A2(new_n672), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n618), .A2(new_n672), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n630), .A2(new_n633), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n687), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n630), .B1(new_n939), .B2(new_n525), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n942), .A2(KEYINPUT42), .B1(new_n673), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n541), .A2(new_n672), .ZN(new_n946));
  MUX2_X1   g0746(.A(new_n646), .B(new_n702), .S(new_n946), .Z(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT105), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n943), .A2(new_n945), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n685), .A2(new_n940), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n692), .B(new_n954), .Z(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n689), .A2(new_n940), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT45), .Z(new_n958));
  NOR2_X1   g0758(.A1(new_n689), .A2(new_n940), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n686), .ZN(new_n962));
  INV_X1    g0762(.A(new_n650), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n684), .B1(new_n963), .B2(new_n672), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(new_n687), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n965), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n965), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n732), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n962), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n956), .B1(new_n973), .B2(new_n733), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n953), .B1(new_n974), .B2(new_n738), .ZN(new_n975));
  INV_X1    g0775(.A(new_n808), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n801), .B1(new_n210), .B2(new_n359), .C1(new_n976), .C2(new_n235), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n977), .A2(new_n739), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n281), .B1(new_n780), .B2(new_n785), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G58), .B2(new_n788), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n769), .A2(G150), .B1(new_n750), .B2(G143), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G50), .A2(new_n782), .B1(new_n777), .B2(G137), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n755), .A2(new_n324), .ZN(new_n983));
  INV_X1    g0783(.A(new_n758), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(G77), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n756), .A2(new_n509), .B1(new_n984), .B2(G97), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G283), .A2(new_n782), .B1(new_n777), .B2(G317), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n463), .A3(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n472), .A2(new_n764), .B1(new_n769), .B2(G303), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n745), .B2(new_n588), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  XOR2_X1   g0793(.A(KEYINPUT108), .B(G311), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n750), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n986), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n978), .B1(new_n743), .B2(new_n998), .C1(new_n948), .C2(new_n813), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n975), .A2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n684), .A2(new_n800), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n694), .A2(new_n803), .B1(G107), .B2(new_n210), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n694), .B(new_n479), .C1(new_n324), .C2(new_n328), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT109), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n258), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n1006), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT50), .B1(new_n1006), .B2(G50), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n976), .B1(new_n232), .B2(G45), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1002), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT110), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n801), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n739), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n761), .A2(new_n533), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n258), .A2(new_n764), .B1(new_n750), .B2(G159), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n324), .B2(new_n773), .ZN(new_n1018));
  XOR2_X1   g0818(.A(KEYINPUT111), .B(G150), .Z(new_n1019));
  OAI221_X1 g0819(.A(new_n394), .B1(new_n776), .B2(new_n1019), .C1(new_n770), .C2(new_n202), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n755), .A2(new_n359), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n745), .A2(new_n328), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR4_X1    g0823(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n756), .A2(G283), .B1(new_n788), .B2(new_n472), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n994), .A2(new_n764), .B1(new_n750), .B2(G322), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n769), .A2(G317), .B1(G303), .B2(new_n782), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1025), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n394), .B1(G326), .B2(new_n777), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n588), .C2(new_n758), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1024), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1015), .B1(new_n1037), .B2(new_n742), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n970), .A2(new_n738), .B1(new_n1001), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n692), .B1(new_n971), .B2(new_n732), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n733), .A2(new_n970), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(G393));
  NAND2_X1  g0842(.A1(new_n941), .A2(new_n800), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n394), .B1(new_n819), .B2(new_n776), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1044), .B(new_n831), .C1(G68), .C2(new_n788), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n756), .A2(G77), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n1006), .B2(new_n773), .C1(new_n780), .C2(new_n202), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1047), .A2(KEYINPUT113), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n769), .A2(G159), .B1(new_n750), .B2(G150), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(KEYINPUT113), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n780), .A2(new_n746), .B1(new_n776), .B2(new_n771), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n281), .B(new_n1053), .C1(G294), .C2(new_n782), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n769), .A2(G311), .B1(new_n750), .B2(G317), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n756), .A2(G116), .B1(new_n788), .B2(G283), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1054), .A2(new_n1056), .A3(new_n784), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n743), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n240), .A2(new_n808), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n802), .B1(G97), .B2(new_n691), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n811), .B(new_n1059), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT114), .Z(new_n1063));
  AOI22_X1  g0863(.A1(new_n962), .A2(new_n738), .B1(new_n1043), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n973), .A2(new_n692), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n962), .A2(new_n972), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(G390));
  AND4_X1   g0867(.A1(G330), .A2(new_n917), .A3(new_n844), .A4(new_n910), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n901), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n900), .A2(new_n904), .B1(new_n1069), .B2(new_n911), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n839), .B1(new_n707), .B2(new_n838), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n910), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n916), .A2(new_n901), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1068), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n911), .A2(new_n1069), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n891), .B1(new_n890), .B2(new_n899), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n903), .A2(KEYINPUT103), .A3(new_n898), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n730), .A2(new_n844), .A3(new_n910), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1082), .A3(new_n1075), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n738), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n799), .B1(new_n900), .B2(new_n904), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n769), .A2(G132), .B1(G125), .B2(new_n777), .ZN(new_n1087));
  INV_X1    g0887(.A(G128), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT119), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1087), .B1(new_n1088), .B2(new_n751), .C1(new_n1091), .C2(new_n773), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n409), .B1(new_n764), .B2(G137), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n202), .B2(new_n758), .C1(new_n785), .C2(new_n755), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1019), .A2(new_n745), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT53), .Z(new_n1096));
  NOR3_X1   g0896(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n761), .A2(new_n324), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n780), .A2(new_n351), .B1(new_n751), .B2(new_n825), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n281), .B1(new_n777), .B2(G294), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1046), .B(new_n1100), .C1(new_n512), .C2(new_n745), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n770), .A2(new_n588), .B1(new_n773), .B2(new_n533), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n742), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1104), .B(new_n739), .C1(new_n258), .C2(new_n835), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1086), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT120), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1085), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n462), .A2(new_n730), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n851), .A2(new_n665), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n839), .B1(new_n699), .B2(new_n844), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n917), .A2(G330), .A3(new_n844), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1072), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1113), .B1(new_n1115), .B2(new_n1082), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT115), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n910), .B1(new_n730), .B2(new_n844), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1068), .A2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1116), .A2(new_n1117), .B1(new_n1119), .B2(new_n1071), .ZN(new_n1120));
  OAI21_X1  g0920(.A(KEYINPUT115), .B1(new_n1119), .B2(new_n1113), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1112), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1077), .A2(new_n1083), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT116), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1077), .A2(new_n1083), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(KEYINPUT117), .A3(new_n692), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1084), .A2(new_n1122), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n693), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT118), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1129), .B1(new_n1132), .B2(KEYINPUT117), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT118), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1110), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G378));
  NAND2_X1  g0940(.A1(new_n921), .A2(G330), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT121), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n265), .A2(new_n670), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n664), .A2(new_n345), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n345), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n302), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  NAND3_X1  g0950(.A1(new_n1145), .A2(new_n1147), .A3(new_n1142), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1141), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n921), .B(G330), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT122), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(new_n912), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n738), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n739), .B1(G50), .B2(new_n835), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n394), .A2(G41), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G50), .B(new_n1161), .C1(new_n268), .C2(new_n269), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n770), .A2(new_n493), .B1(new_n776), .B2(new_n825), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n758), .A2(new_n371), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1163), .A2(new_n983), .A3(new_n1022), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n764), .A2(G97), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n750), .A2(G116), .B1(new_n567), .B2(new_n782), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1165), .A2(new_n1161), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT58), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(G132), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n780), .A2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n770), .A2(new_n1088), .B1(new_n773), .B2(new_n818), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G125), .C2(new_n750), .ZN(new_n1174));
  INV_X1    g0974(.A(G150), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n755), .C1(new_n745), .C2(new_n1091), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n984), .A2(G159), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1170), .B1(new_n1169), .B2(new_n1168), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1160), .B1(new_n1182), .B2(new_n742), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1154), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n799), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1112), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1127), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1158), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1112), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n912), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n912), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n692), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1159), .B(new_n1185), .C1(new_n1188), .C2(new_n1194), .ZN(G375));
  INV_X1    g0995(.A(new_n1122), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1120), .A2(new_n1112), .A3(new_n1121), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n955), .A3(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT123), .Z(new_n1199));
  AOI21_X1  g0999(.A(new_n737), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1072), .A2(new_n798), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n739), .B1(G68), .B2(new_n835), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n770), .A2(new_n818), .B1(new_n751), .B2(new_n1171), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n773), .A2(new_n1175), .B1(new_n776), .B2(new_n1088), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1090), .A2(new_n764), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1164), .A2(new_n463), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n756), .A2(G50), .B1(new_n788), .B2(G159), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n588), .A2(new_n780), .B1(new_n770), .B2(new_n825), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G294), .B2(new_n750), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n773), .A2(new_n351), .B1(new_n776), .B2(new_n746), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1021), .B(new_n1212), .C1(G97), .C2(new_n788), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n409), .B1(new_n761), .B2(new_n328), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1211), .B(new_n1213), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1215), .A2(new_n1214), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1209), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1202), .B1(new_n1218), .B2(new_n742), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1200), .B1(new_n1201), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1199), .A2(new_n1220), .ZN(G381));
  OR2_X1    g1021(.A1(G393), .A2(G396), .ZN(new_n1222));
  OR4_X1    g1022(.A1(G384), .A2(G387), .A3(new_n1222), .A4(G390), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1110), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G375), .A2(new_n1223), .A3(G381), .A4(new_n1225), .ZN(G407));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1227), .A2(G213), .A3(new_n671), .A4(new_n1224), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G407), .A2(G213), .A3(new_n1228), .ZN(G409));
  XNOR2_X1  g1029(.A(G387), .B(G390), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(G393), .B(new_n815), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1230), .B(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n671), .A2(G213), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1196), .A2(KEYINPUT60), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1234), .A2(new_n1197), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n692), .B1(new_n1234), .B2(new_n1197), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1220), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(new_n849), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n849), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G375), .B1(new_n1241), .B2(new_n1109), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n738), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1185), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1187), .A2(new_n1158), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n955), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1225), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1233), .B(new_n1240), .C1(new_n1242), .C2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1139), .A2(G375), .B1(new_n1225), .B2(new_n1246), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1251), .A2(KEYINPUT125), .A3(new_n1233), .A4(new_n1240), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT62), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1254));
  OAI21_X1  g1054(.A(new_n1233), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1240), .B(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1248), .A2(KEYINPUT62), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1232), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1250), .A2(new_n1252), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1233), .A4(new_n1240), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1232), .A2(KEYINPUT61), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1261), .A2(new_n1267), .ZN(G405));
  INV_X1    g1068(.A(new_n1242), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G375), .A2(new_n1224), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1240), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1240), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1273), .A3(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(new_n1232), .ZN(G402));
endmodule


