

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U559 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n543) );
  NOR2_X2 U560 ( .A1(G164), .A2(G1384), .ZN(n716) );
  XOR2_X1 U561 ( .A(n729), .B(KEYINPUT92), .Z(n726) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n723) );
  XOR2_X1 U563 ( .A(n566), .B(KEYINPUT66), .Z(n524) );
  XOR2_X1 U564 ( .A(KEYINPUT79), .B(n533), .Z(n525) );
  NOR2_X1 U565 ( .A1(n740), .A2(n739), .ZN(n741) );
  INV_X1 U566 ( .A(KEYINPUT31), .ZN(n764) );
  NOR2_X1 U567 ( .A1(n797), .A2(n796), .ZN(n803) );
  XOR2_X1 U568 ( .A(KEYINPUT15), .B(n602), .Z(n987) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  XNOR2_X1 U570 ( .A(KEYINPUT80), .B(n541), .ZN(G168) );
  INV_X1 U571 ( .A(G651), .ZN(n534) );
  NOR2_X1 U572 ( .A1(n640), .A2(n534), .ZN(n650) );
  NAND2_X1 U573 ( .A1(G76), .A2(n650), .ZN(n529) );
  XOR2_X1 U574 ( .A(KEYINPUT77), .B(KEYINPUT4), .Z(n527) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U576 ( .A1(G89), .A2(n654), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n530), .B(KEYINPUT78), .ZN(n531) );
  XNOR2_X1 U580 ( .A(KEYINPUT5), .B(n531), .ZN(n539) );
  NOR2_X1 U581 ( .A1(G651), .A2(n640), .ZN(n532) );
  XNOR2_X2 U582 ( .A(KEYINPUT64), .B(n532), .ZN(n659) );
  NAND2_X1 U583 ( .A1(G51), .A2(n659), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X2 U585 ( .A(KEYINPUT1), .B(n535), .Z(n653) );
  NAND2_X1 U586 ( .A1(n653), .A2(G63), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n525), .A2(n536), .ZN(n537) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(n537), .Z(n538) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U590 ( .A(n540), .B(KEYINPUT7), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U592 ( .A(G2105), .ZN(n561) );
  AND2_X1 U593 ( .A1(n561), .A2(G2104), .ZN(n888) );
  NAND2_X1 U594 ( .A1(G102), .A2(n888), .ZN(n545) );
  NOR2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  XNOR2_X2 U596 ( .A(n543), .B(n542), .ZN(n889) );
  NAND2_X1 U597 ( .A1(G138), .A2(n889), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n549) );
  AND2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U600 ( .A1(G114), .A2(n884), .ZN(n547) );
  NOR2_X2 U601 ( .A1(G2104), .A2(n561), .ZN(n885) );
  NAND2_X1 U602 ( .A1(G126), .A2(n885), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n549), .A2(n548), .ZN(G164) );
  NAND2_X1 U605 ( .A1(n653), .A2(G64), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT69), .B(n550), .Z(n552) );
  NAND2_X1 U607 ( .A1(G52), .A2(n659), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U609 ( .A(KEYINPUT70), .B(n553), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G77), .A2(n650), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G90), .A2(n654), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U613 ( .A(KEYINPUT9), .B(n556), .ZN(n557) );
  XNOR2_X1 U614 ( .A(KEYINPUT71), .B(n557), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n559), .A2(n558), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  AND2_X1 U617 ( .A1(G2104), .A2(G101), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT65), .ZN(n563) );
  XNOR2_X1 U620 ( .A(n563), .B(KEYINPUT23), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G125), .A2(n885), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G137), .A2(n889), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G113), .A2(n884), .ZN(n567) );
  AND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n686) );
  AND2_X1 U626 ( .A1(n524), .A2(n686), .ZN(G160) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  NAND2_X1 U630 ( .A1(G75), .A2(n650), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G88), .A2(n654), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G62), .A2(n653), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G50), .A2(n659), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(G166) );
  NAND2_X1 U637 ( .A1(G65), .A2(n653), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G91), .A2(n654), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n650), .A2(G78), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT72), .B(n577), .Z(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G53), .A2(n659), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(G299) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n831) );
  NAND2_X1 U648 ( .A1(n831), .A2(G567), .ZN(n583) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  NAND2_X1 U650 ( .A1(G56), .A2(n653), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n584), .Z(n591) );
  NAND2_X1 U652 ( .A1(G81), .A2(n654), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT12), .ZN(n586) );
  XNOR2_X1 U654 ( .A(n586), .B(KEYINPUT74), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G68), .A2(n650), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U657 ( .A(KEYINPUT13), .B(n589), .Z(n590) );
  NOR2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U659 ( .A1(G43), .A2(n659), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n982) );
  INV_X1 U661 ( .A(G860), .ZN(n629) );
  OR2_X1 U662 ( .A1(n982), .A2(n629), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G92), .A2(n654), .ZN(n594) );
  XNOR2_X1 U665 ( .A(n594), .B(KEYINPUT76), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G79), .A2(n650), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G54), .A2(n659), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G66), .A2(n653), .ZN(n597) );
  XNOR2_X1 U670 ( .A(KEYINPUT75), .B(n597), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  INV_X1 U673 ( .A(G868), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n987), .A2(n605), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G284) );
  NOR2_X1 U676 ( .A1(G286), .A2(n605), .ZN(n606) );
  XOR2_X1 U677 ( .A(KEYINPUT81), .B(n606), .Z(n608) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n629), .A2(G559), .ZN(n609) );
  INV_X1 U681 ( .A(n987), .ZN(n626) );
  NAND2_X1 U682 ( .A1(n609), .A2(n626), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT82), .ZN(n611) );
  XNOR2_X1 U684 ( .A(KEYINPUT16), .B(n611), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n982), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G868), .A2(n626), .ZN(n612) );
  NOR2_X1 U687 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G99), .A2(n888), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G111), .A2(n884), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U692 ( .A(KEYINPUT84), .B(n617), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G123), .A2(n885), .ZN(n618) );
  XOR2_X1 U694 ( .A(KEYINPUT18), .B(n618), .Z(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(KEYINPUT83), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G135), .A2(n889), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n949) );
  XNOR2_X1 U699 ( .A(n949), .B(G2096), .ZN(n625) );
  INV_X1 U700 ( .A(G2100), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(G156) );
  XNOR2_X1 U702 ( .A(n982), .B(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n626), .A2(G559), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n628), .B(n627), .ZN(n667) );
  NAND2_X1 U705 ( .A1(n629), .A2(n667), .ZN(n636) );
  NAND2_X1 U706 ( .A1(G67), .A2(n653), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G55), .A2(n659), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G80), .A2(n650), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G93), .A2(n654), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n669) );
  XOR2_X1 U713 ( .A(n636), .B(n669), .Z(G145) );
  NAND2_X1 U714 ( .A1(G651), .A2(G74), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G49), .A2(n659), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U717 ( .A1(n653), .A2(n639), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n640), .A2(G87), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G85), .A2(n654), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G47), .A2(n659), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G72), .A2(n650), .ZN(n645) );
  XOR2_X1 U724 ( .A(KEYINPUT68), .B(n645), .Z(n646) );
  NOR2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n653), .A2(G60), .ZN(n648) );
  NAND2_X1 U727 ( .A1(n649), .A2(n648), .ZN(G290) );
  XOR2_X1 U728 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n652) );
  NAND2_X1 U729 ( .A1(G73), .A2(n650), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n652), .B(n651), .ZN(n658) );
  NAND2_X1 U731 ( .A1(G61), .A2(n653), .ZN(n656) );
  NAND2_X1 U732 ( .A1(G86), .A2(n654), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U735 ( .A1(G48), .A2(n659), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n661), .A2(n660), .ZN(G305) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(G288), .ZN(n666) );
  XNOR2_X1 U738 ( .A(G166), .B(n669), .ZN(n664) );
  XNOR2_X1 U739 ( .A(G290), .B(G299), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(G305), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n666), .B(n665), .ZN(n902) );
  XNOR2_X1 U743 ( .A(n667), .B(n902), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n668), .A2(G868), .ZN(n671) );
  OR2_X1 U745 ( .A1(G868), .A2(n669), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n671), .A2(n670), .ZN(G295) );
  INV_X1 U747 ( .A(G2072), .ZN(n945) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT21), .B(n674), .Z(n675) );
  NOR2_X1 U752 ( .A1(n945), .A2(n675), .ZN(n676) );
  XNOR2_X1 U753 ( .A(KEYINPUT87), .B(n676), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U755 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U756 ( .A1(G219), .A2(G220), .ZN(n677) );
  XOR2_X1 U757 ( .A(KEYINPUT88), .B(n677), .Z(n678) );
  XNOR2_X1 U758 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  NOR2_X1 U759 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G96), .A2(n680), .ZN(n836) );
  NAND2_X1 U761 ( .A1(n836), .A2(G2106), .ZN(n684) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n681) );
  NOR2_X1 U763 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U764 ( .A1(G108), .A2(n682), .ZN(n837) );
  NAND2_X1 U765 ( .A1(n837), .A2(G567), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n858) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n858), .A2(n685), .ZN(n835) );
  NAND2_X1 U769 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U771 ( .A(G1986), .B(G290), .ZN(n984) );
  AND2_X1 U772 ( .A1(G40), .A2(n686), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n687), .A2(n524), .ZN(n717) );
  NOR2_X1 U774 ( .A1(n716), .A2(n717), .ZN(n826) );
  NAND2_X1 U775 ( .A1(n984), .A2(n826), .ZN(n815) );
  XNOR2_X1 U776 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NAND2_X1 U777 ( .A1(n889), .A2(G140), .ZN(n688) );
  XOR2_X1 U778 ( .A(KEYINPUT89), .B(n688), .Z(n690) );
  NAND2_X1 U779 ( .A1(n888), .A2(G104), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U781 ( .A(KEYINPUT34), .B(n691), .ZN(n696) );
  NAND2_X1 U782 ( .A1(G116), .A2(n884), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G128), .A2(n885), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U785 ( .A(KEYINPUT35), .B(n694), .Z(n695) );
  NOR2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U787 ( .A(KEYINPUT36), .B(n697), .ZN(n899) );
  NOR2_X1 U788 ( .A1(n824), .A2(n899), .ZN(n964) );
  NAND2_X1 U789 ( .A1(n826), .A2(n964), .ZN(n822) );
  NAND2_X1 U790 ( .A1(G117), .A2(n884), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G129), .A2(n885), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n888), .A2(G105), .ZN(n700) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n700), .Z(n701) );
  NOR2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n889), .A2(G141), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n867) );
  NAND2_X1 U798 ( .A1(G1996), .A2(n867), .ZN(n705) );
  XNOR2_X1 U799 ( .A(n705), .B(KEYINPUT90), .ZN(n713) );
  NAND2_X1 U800 ( .A1(G95), .A2(n888), .ZN(n707) );
  NAND2_X1 U801 ( .A1(G107), .A2(n884), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U803 ( .A1(G131), .A2(n889), .ZN(n709) );
  NAND2_X1 U804 ( .A1(G119), .A2(n885), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n868) );
  NAND2_X1 U807 ( .A1(G1991), .A2(n868), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n960) );
  NAND2_X1 U809 ( .A1(n960), .A2(n826), .ZN(n714) );
  XNOR2_X1 U810 ( .A(n714), .B(KEYINPUT91), .ZN(n819) );
  INV_X1 U811 ( .A(n819), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n822), .A2(n715), .ZN(n813) );
  INV_X1 U813 ( .A(n716), .ZN(n718) );
  NOR2_X2 U814 ( .A1(n718), .A2(n717), .ZN(n729) );
  NOR2_X1 U815 ( .A1(n726), .A2(n945), .ZN(n720) );
  XNOR2_X1 U816 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n719) );
  XNOR2_X1 U817 ( .A(n720), .B(n719), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n726), .A2(G1956), .ZN(n743) );
  INV_X1 U819 ( .A(G299), .ZN(n721) );
  AND2_X1 U820 ( .A1(n743), .A2(n721), .ZN(n722) );
  NAND2_X1 U821 ( .A1(n744), .A2(n722), .ZN(n724) );
  XNOR2_X1 U822 ( .A(n724), .B(n723), .ZN(n742) );
  INV_X1 U823 ( .A(n729), .ZN(n769) );
  NAND2_X1 U824 ( .A1(G1348), .A2(n769), .ZN(n725) );
  XNOR2_X1 U825 ( .A(n725), .B(KEYINPUT96), .ZN(n728) );
  INV_X1 U826 ( .A(n726), .ZN(n751) );
  NAND2_X1 U827 ( .A1(G2067), .A2(n751), .ZN(n727) );
  NAND2_X1 U828 ( .A1(n728), .A2(n727), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n738), .A2(n987), .ZN(n737) );
  INV_X1 U830 ( .A(n982), .ZN(n735) );
  NAND2_X1 U831 ( .A1(G1996), .A2(n729), .ZN(n730) );
  XNOR2_X1 U832 ( .A(n730), .B(KEYINPUT26), .ZN(n732) );
  NAND2_X1 U833 ( .A1(G1341), .A2(n769), .ZN(n731) );
  NAND2_X1 U834 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U835 ( .A(n733), .B(KEYINPUT95), .ZN(n734) );
  AND2_X1 U836 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n740) );
  NOR2_X1 U838 ( .A1(n987), .A2(n738), .ZN(n739) );
  NAND2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U841 ( .A1(G299), .A2(n745), .ZN(n746) );
  XNOR2_X1 U842 ( .A(n746), .B(KEYINPUT28), .ZN(n747) );
  NAND2_X1 U843 ( .A1(n748), .A2(n747), .ZN(n750) );
  XNOR2_X1 U844 ( .A(KEYINPUT98), .B(KEYINPUT29), .ZN(n749) );
  XNOR2_X1 U845 ( .A(n750), .B(n749), .ZN(n756) );
  XNOR2_X1 U846 ( .A(G2078), .B(KEYINPUT25), .ZN(n936) );
  NAND2_X1 U847 ( .A1(n751), .A2(n936), .ZN(n753) );
  INV_X1 U848 ( .A(G1961), .ZN(n1006) );
  NAND2_X1 U849 ( .A1(n769), .A2(n1006), .ZN(n752) );
  NAND2_X1 U850 ( .A1(n753), .A2(n752), .ZN(n761) );
  AND2_X1 U851 ( .A1(n761), .A2(G171), .ZN(n754) );
  XOR2_X1 U852 ( .A(KEYINPUT93), .B(n754), .Z(n755) );
  NOR2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U854 ( .A(KEYINPUT99), .B(n757), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n769), .A2(G8), .ZN(n796) );
  NOR2_X1 U856 ( .A1(G1966), .A2(n796), .ZN(n782) );
  NOR2_X1 U857 ( .A1(G2084), .A2(n769), .ZN(n778) );
  NOR2_X1 U858 ( .A1(n782), .A2(n778), .ZN(n758) );
  NAND2_X1 U859 ( .A1(G8), .A2(n758), .ZN(n759) );
  XNOR2_X1 U860 ( .A(KEYINPUT30), .B(n759), .ZN(n760) );
  NOR2_X1 U861 ( .A1(G168), .A2(n760), .ZN(n763) );
  NOR2_X1 U862 ( .A1(G171), .A2(n761), .ZN(n762) );
  NOR2_X1 U863 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U864 ( .A(n765), .B(n764), .ZN(n766) );
  NAND2_X1 U865 ( .A1(n767), .A2(n766), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n780), .A2(G286), .ZN(n768) );
  XNOR2_X1 U867 ( .A(n768), .B(KEYINPUT100), .ZN(n775) );
  NOR2_X1 U868 ( .A1(G1971), .A2(n796), .ZN(n771) );
  NOR2_X1 U869 ( .A1(G2090), .A2(n769), .ZN(n770) );
  NOR2_X1 U870 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U871 ( .A1(n772), .A2(G303), .ZN(n773) );
  XOR2_X1 U872 ( .A(KEYINPUT101), .B(n773), .Z(n774) );
  NAND2_X1 U873 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n776), .A2(G8), .ZN(n777) );
  XOR2_X1 U875 ( .A(KEYINPUT32), .B(n777), .Z(n784) );
  NAND2_X1 U876 ( .A1(G8), .A2(n778), .ZN(n779) );
  NAND2_X1 U877 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U878 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X2 U879 ( .A1(n784), .A2(n783), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G166), .A2(G8), .ZN(n785) );
  NOR2_X1 U881 ( .A1(G2090), .A2(n785), .ZN(n786) );
  NOR2_X1 U882 ( .A1(n795), .A2(n786), .ZN(n787) );
  XNOR2_X1 U883 ( .A(KEYINPUT103), .B(n787), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n788), .A2(n796), .ZN(n792) );
  INV_X1 U885 ( .A(n796), .ZN(n799) );
  NOR2_X1 U886 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XNOR2_X1 U887 ( .A(n789), .B(KEYINPUT24), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n799), .A2(n790), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n811) );
  XNOR2_X1 U890 ( .A(G1981), .B(G305), .ZN(n972) );
  NOR2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n798) );
  INV_X1 U892 ( .A(n798), .ZN(n794) );
  INV_X1 U893 ( .A(G1971), .ZN(n974) );
  NAND2_X1 U894 ( .A1(G166), .A2(n974), .ZN(n793) );
  NAND2_X1 U895 ( .A1(n794), .A2(n793), .ZN(n976) );
  NOR2_X1 U896 ( .A1(n795), .A2(n976), .ZN(n797) );
  NAND2_X1 U897 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U898 ( .A(KEYINPUT33), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U900 ( .A1(n805), .A2(n800), .ZN(n801) );
  XOR2_X1 U901 ( .A(n801), .B(KEYINPUT102), .Z(n804) );
  AND2_X1 U902 ( .A1(n977), .A2(n804), .ZN(n802) );
  NAND2_X1 U903 ( .A1(n803), .A2(n802), .ZN(n808) );
  INV_X1 U904 ( .A(n804), .ZN(n806) );
  OR2_X1 U905 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n972), .A2(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n829) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n867), .ZN(n952) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n868), .ZN(n950) );
  NOR2_X1 U914 ( .A1(n816), .A2(n950), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n817), .B(KEYINPUT104), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n952), .A2(n820), .ZN(n821) );
  XNOR2_X1 U918 ( .A(KEYINPUT39), .B(n821), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n824), .A2(n899), .ZN(n965) );
  NAND2_X1 U921 ( .A1(n825), .A2(n965), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n832) );
  XNOR2_X1 U927 ( .A(KEYINPUT107), .B(n832), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n833), .A2(G661), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U936 ( .A(G1996), .B(KEYINPUT41), .ZN(n847) );
  XOR2_X1 U937 ( .A(G1981), .B(G1956), .Z(n839) );
  XNOR2_X1 U938 ( .A(G1991), .B(G1966), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1961), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(G2474), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U948 ( .A(KEYINPUT108), .B(G2678), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2090), .Z(n851) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U953 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U954 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G227) );
  INV_X1 U958 ( .A(n858), .ZN(G319) );
  NAND2_X1 U959 ( .A1(G124), .A2(n885), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n859), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G136), .A2(n889), .ZN(n860) );
  XOR2_X1 U962 ( .A(KEYINPUT111), .B(n860), .Z(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G100), .A2(n888), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G112), .A2(n884), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U967 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U968 ( .A(G164), .B(n867), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n871) );
  XNOR2_X1 U971 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n883) );
  NAND2_X1 U974 ( .A1(G103), .A2(n888), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G139), .A2(n889), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n884), .A2(G115), .ZN(n876) );
  XOR2_X1 U978 ( .A(KEYINPUT113), .B(n876), .Z(n878) );
  NAND2_X1 U979 ( .A1(n885), .A2(G127), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n944) );
  XNOR2_X1 U983 ( .A(G160), .B(n944), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n896) );
  NAND2_X1 U985 ( .A1(G118), .A2(n884), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G130), .A2(n885), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U988 ( .A1(G106), .A2(n888), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U991 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U993 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U994 ( .A(G162), .B(n949), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n900) );
  XOR2_X1 U996 ( .A(n900), .B(n899), .Z(n901) );
  NOR2_X1 U997 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U998 ( .A(n902), .B(G286), .ZN(n905) );
  XOR2_X1 U999 ( .A(KEYINPUT115), .B(n982), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n987), .B(n903), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(G301), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n922) );
  XNOR2_X1 U1007 ( .A(G2454), .B(G2427), .ZN(n919) );
  XOR2_X1 U1008 ( .A(KEYINPUT106), .B(G2430), .Z(n911) );
  XNOR2_X1 U1009 ( .A(G2443), .B(G2451), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1011 ( .A(G2446), .B(KEYINPUT105), .Z(n913) );
  XNOR2_X1 U1012 ( .A(G1348), .B(G1341), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1014 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1015 ( .A(G2435), .B(G2438), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(G14), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n925), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G96), .ZN(G221) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1027 ( .A(G2090), .B(G35), .Z(n928) );
  XOR2_X1 U1028 ( .A(G34), .B(KEYINPUT54), .Z(n926) );
  XNOR2_X1 U1029 ( .A(G2084), .B(n926), .ZN(n927) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(G1991), .B(G25), .ZN(n929) );
  NOR2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G33), .B(n945), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n931), .A2(G28), .ZN(n933) );
  XNOR2_X1 U1036 ( .A(G32), .B(G1996), .ZN(n932) );
  NOR2_X1 U1037 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1039 ( .A(G27), .B(n936), .Z(n937) );
  NOR2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(n939), .B(KEYINPUT53), .ZN(n940) );
  NOR2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(G29), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(n943), .B(KEYINPUT55), .ZN(n970) );
  XOR2_X1 U1045 ( .A(G164), .B(G2078), .Z(n947) );
  XNOR2_X1 U1046 ( .A(n945), .B(n944), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(KEYINPUT50), .B(n948), .ZN(n962) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n958) );
  XOR2_X1 U1050 ( .A(G160), .B(G2084), .Z(n956) );
  XOR2_X1 U1051 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1053 ( .A(KEYINPUT51), .B(n953), .Z(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT117), .B(n954), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(G29), .A2(n968), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n1029) );
  XOR2_X1 U1064 ( .A(G168), .B(G1966), .Z(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT57), .B(n973), .Z(n992) );
  NOR2_X1 U1067 ( .A1(G166), .A2(n974), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G299), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT120), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n987), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT118), .B(n988), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G1961), .B(G301), .Z(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT119), .B(n993), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1083 ( .A(KEYINPUT56), .B(G16), .Z(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n1025) );
  XOR2_X1 U1085 ( .A(G16), .B(KEYINPUT121), .Z(n1023) );
  XNOR2_X1 U1086 ( .A(G1986), .B(G24), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT122), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT123), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT124), .ZN(n1020) );
  XOR2_X1 U1095 ( .A(G1966), .B(G21), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G5), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1018) );
  XOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT59), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G20), .B(G1956), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G1341), .B(G19), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G1981), .B(G6), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT60), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(n1021), .B(KEYINPUT61), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT125), .B(n1026), .Z(n1027) );
  NAND2_X1 U1113 ( .A1(G11), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(n1031), .B(n1030), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
endmodule

