//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT17), .ZN(new_n189));
  INV_X1    g003(.A(G131), .ZN(new_n190));
  NOR2_X1   g004(.A1(G237), .A2(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(G214), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT91), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT91), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G214), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(new_n194), .ZN(new_n198));
  AOI211_X1 g012(.A(new_n189), .B(new_n190), .C1(new_n196), .C2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n202), .B1(new_n206), .B2(new_n200), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(G146), .B(new_n202), .C1(new_n206), .C2(new_n200), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT94), .B1(new_n199), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n190), .B1(new_n196), .B2(new_n198), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT17), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT94), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n209), .A4(new_n210), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n197), .B1(new_n193), .B2(new_n194), .ZN(new_n217));
  INV_X1    g031(.A(new_n198), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n196), .A2(new_n190), .A3(new_n198), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n189), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n212), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G125), .B(G140), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(new_n208), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n196), .A2(new_n198), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(new_n190), .ZN(new_n227));
  OAI221_X1 g041(.A(new_n224), .B1(new_n225), .B2(new_n227), .C1(new_n219), .C2(new_n226), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT93), .B(G104), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n229), .B(new_n230), .Z(new_n231));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n196), .A2(new_n190), .A3(new_n198), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT92), .B1(new_n233), .B2(new_n213), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(new_n235), .A3(new_n220), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT19), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n206), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n223), .A2(KEYINPUT19), .ZN(new_n239));
  AOI21_X1  g053(.A(G146), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n210), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n228), .ZN(new_n244));
  INV_X1    g058(.A(new_n231), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT20), .B(new_n188), .C1(new_n232), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n232), .A2(new_n246), .A3(KEYINPUT95), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT95), .B1(new_n232), .B2(new_n246), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n249), .A2(new_n250), .A3(new_n188), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  AOI211_X1 g069(.A(new_n254), .B(new_n255), .C1(G234), .C2(G237), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT21), .B(G898), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(G234), .A2(G237), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT99), .A2(G952), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT99), .A2(G952), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n255), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n222), .A2(new_n228), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n245), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n232), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n254), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G475), .ZN(new_n269));
  XNOR2_X1  g083(.A(G128), .B(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n272), .A2(KEYINPUT13), .A3(G143), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n274), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT97), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n271), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G107), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT96), .B1(new_n280), .B2(G122), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT96), .ZN(new_n282));
  INV_X1    g096(.A(G122), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(G122), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n279), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(new_n279), .A3(new_n286), .ZN(new_n288));
  OAI221_X1 g102(.A(new_n278), .B1(new_n277), .B2(new_n276), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n281), .A2(new_n284), .B1(new_n286), .B2(KEYINPUT14), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n290), .A2(KEYINPUT98), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n290), .B2(KEYINPUT98), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n279), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n270), .B(G134), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n295), .A2(new_n288), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n289), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  INV_X1    g112(.A(G217), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(new_n299), .A3(G953), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n301), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G478), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT15), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n253), .A2(new_n264), .A3(new_n269), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT100), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n232), .A2(new_n246), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n232), .A2(new_n246), .A3(KEYINPUT95), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n187), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n247), .B1(new_n314), .B2(KEYINPUT20), .ZN(new_n315));
  INV_X1    g129(.A(new_n269), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT100), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n264), .A4(new_n307), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n309), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G122), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT85), .A2(KEYINPUT6), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n279), .A3(G104), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n324), .A2(new_n327), .A3(new_n279), .A4(G104), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n279), .A2(G104), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT80), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n326), .A2(new_n334), .A3(new_n328), .A4(new_n330), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n333), .A3(G101), .A4(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT2), .B(G113), .Z(new_n337));
  XNOR2_X1  g151(.A(G116), .B(G119), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n337), .A2(KEYINPUT69), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT69), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n339), .A2(new_n340), .B1(new_n338), .B2(new_n337), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n332), .A2(G101), .A3(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(G101), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n326), .A2(new_n344), .A3(new_n328), .A4(new_n330), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n343), .A2(KEYINPUT81), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT81), .B1(new_n343), .B2(new_n346), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G107), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n351), .B2(new_n329), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G119), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G116), .ZN(new_n358));
  OAI21_X1  g172(.A(G113), .B1(new_n358), .B2(KEYINPUT5), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n339), .A2(new_n340), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(new_n322), .B(new_n323), .C1(new_n349), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n322), .B1(new_n349), .B2(new_n362), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n349), .A2(new_n362), .A3(new_n322), .ZN(new_n366));
  INV_X1    g180(.A(new_n323), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n363), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n208), .A2(G143), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n371));
  INV_X1    g185(.A(G143), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G146), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n371), .B1(new_n372), .B2(G146), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OR3_X1    g190(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n377), .A2(new_n378), .B1(KEYINPUT0), .B2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(G146), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n370), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT0), .A3(G128), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n204), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT1), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n388), .A3(G128), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n372), .C2(G146), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G128), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT67), .B1(new_n370), .B2(KEYINPUT1), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(KEYINPUT65), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n394), .A2(new_n373), .B1(G143), .B2(new_n208), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT68), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT1), .B1(new_n372), .B2(G146), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT67), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(G128), .A3(new_n390), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT68), .B1(new_n401), .B2(new_n376), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n389), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n387), .B1(new_n403), .B2(G125), .ZN(new_n404));
  INV_X1    g218(.A(new_n389), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n396), .B1(new_n393), .B2(new_n395), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n376), .A3(KEYINPUT68), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT86), .A3(new_n204), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n386), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G224), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G953), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n321), .B1(new_n369), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n412), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n410), .B(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(KEYINPUT87), .C1(new_n417), .C2(new_n363), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n415), .A2(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n404), .A2(new_n409), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n386), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n404), .A2(KEYINPUT89), .A3(new_n409), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n410), .A2(new_n421), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n360), .A2(new_n353), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n322), .B(KEYINPUT8), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n339), .A2(new_n340), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n356), .A2(KEYINPUT88), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n359), .B1(new_n355), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n428), .B(new_n429), .C1(new_n354), .C2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n366), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n254), .B1(new_n426), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n419), .A2(new_n420), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n420), .B(KEYINPUT90), .Z(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n414), .B2(new_n418), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n320), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G472), .A2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT32), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n449));
  OR2_X1    g263(.A1(KEYINPUT66), .A2(G137), .ZN(new_n450));
  NAND2_X1  g264(.A1(KEYINPUT66), .A2(G137), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n274), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G134), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n190), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n450), .A2(KEYINPUT11), .A3(G134), .A4(new_n451), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT11), .B1(new_n454), .B2(G134), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n455), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n457), .A2(new_n459), .A3(new_n190), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n403), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n190), .B1(new_n457), .B2(new_n459), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n380), .B(new_n383), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n449), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n461), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n449), .B(new_n464), .C1(new_n408), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n341), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n341), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n462), .A2(new_n470), .A3(new_n464), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT26), .B(G101), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n191), .A2(G210), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n471), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n464), .B1(new_n408), .B2(new_n466), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT30), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n467), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n484), .B2(new_n341), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT71), .A3(new_n477), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT31), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n470), .B1(new_n483), .B2(new_n467), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n489), .A2(new_n481), .A3(new_n476), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n471), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n482), .B(new_n470), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n488), .A2(new_n490), .B1(new_n495), .B2(new_n476), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n487), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n487), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n448), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n476), .B1(new_n489), .B2(new_n481), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(new_n502), .C1(new_n495), .C2(new_n476), .ZN(new_n503));
  MUX2_X1   g317(.A(new_n481), .B(new_n493), .S(KEYINPUT28), .Z(new_n504));
  NOR2_X1   g318(.A1(new_n476), .A2(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n254), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G472), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n487), .A2(new_n496), .A3(new_n497), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n446), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n500), .B(new_n508), .C1(new_n512), .C2(KEYINPUT32), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT77), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n272), .A2(G119), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n357), .A2(G128), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT24), .B(G110), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n515), .B1(KEYINPUT74), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n521), .B(new_n516), .C1(new_n522), .C2(new_n515), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n519), .B1(new_n523), .B2(G110), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n210), .C1(G146), .C2(new_n206), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n517), .A2(new_n518), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n523), .B2(G110), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n211), .A2(new_n527), .A3(KEYINPUT75), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT75), .B1(new_n211), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n525), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT22), .B(G137), .ZN(new_n534));
  INV_X1    g348(.A(G221), .ZN(new_n535));
  INV_X1    g349(.A(G234), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(new_n536), .A3(G953), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n534), .B(new_n537), .Z(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n530), .A2(KEYINPUT76), .A3(new_n538), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n299), .B1(G234), .B2(new_n254), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n542), .B2(new_n543), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n514), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n540), .A2(new_n541), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT25), .B1(new_n549), .B2(G902), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(KEYINPUT77), .A3(new_n544), .A4(new_n546), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n546), .A2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n298), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n535), .B1(new_n559), .B2(new_n254), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n272), .B1(new_n370), .B2(KEYINPUT1), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n389), .B1(new_n382), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n353), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n353), .A2(KEYINPUT10), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n408), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n385), .A2(new_n336), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n348), .B2(new_n347), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n460), .A2(new_n463), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n343), .A2(new_n346), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT81), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n343), .A2(KEYINPUT81), .A3(new_n346), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n570), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(new_n568), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G140), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n255), .A2(G227), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT12), .B1(new_n575), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n353), .A2(new_n563), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n408), .B2(new_n354), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n590), .B2(new_n573), .ZN(new_n591));
  INV_X1    g405(.A(new_n588), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n564), .B1(new_n403), .B2(new_n353), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n575), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n585), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n574), .A3(new_n596), .ZN(new_n597));
  AOI211_X1 g411(.A(G469), .B(G902), .C1(new_n586), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n574), .A2(new_n581), .A3(new_n596), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n580), .A2(new_n568), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(new_n573), .B1(new_n591), .B2(new_n594), .ZN(new_n601));
  OAI211_X1 g415(.A(G469), .B(new_n599), .C1(new_n601), .C2(new_n596), .ZN(new_n602));
  INV_X1    g416(.A(G469), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n254), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n561), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT84), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT84), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n561), .C1(new_n598), .C2(new_n606), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n444), .A2(new_n513), .A3(new_n558), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n614));
  INV_X1    g428(.A(new_n418), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n364), .A2(new_n367), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n578), .A2(new_n579), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n361), .B1(new_n617), .B2(new_n342), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n323), .B1(new_n618), .B2(new_n322), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n364), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT87), .B1(new_n620), .B2(new_n416), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n438), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n420), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n439), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n614), .B1(new_n625), .B2(new_n443), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n420), .B1(new_n419), .B2(new_n438), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n623), .B(new_n437), .C1(new_n414), .C2(new_n418), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n614), .B(new_n443), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n626), .A2(new_n630), .A3(new_n263), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n254), .B1(new_n498), .B2(new_n499), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n445), .B1(new_n498), .B2(new_n499), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n608), .A2(new_n610), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n635), .A2(new_n557), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n302), .A2(new_n303), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT33), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n302), .A2(new_n640), .A3(new_n303), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(G478), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n305), .A2(new_n254), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n304), .B2(new_n305), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n317), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n631), .A2(new_n637), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT102), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  NAND2_X1  g464(.A1(new_n251), .A2(new_n252), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n314), .A2(KEYINPUT20), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n316), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n307), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n631), .A2(new_n637), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT103), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT35), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  AOI21_X1  g474(.A(new_n512), .B1(G472), .B2(new_n632), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n530), .B(new_n662), .Z(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(new_n554), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n548), .A2(new_n551), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n444), .A2(new_n611), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(new_n665), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n510), .A2(new_n511), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n670), .A2(new_n448), .B1(G472), .B2(new_n507), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n634), .A2(new_n447), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n262), .B(KEYINPUT105), .Z(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n256), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT106), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n636), .A2(new_n655), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n443), .B1(new_n627), .B2(new_n628), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n673), .A2(new_n682), .A3(new_n629), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n680), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n611), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT108), .Z(new_n690));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n689), .B(KEYINPUT108), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT109), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n317), .A2(new_n307), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n669), .A2(new_n443), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n442), .B(KEYINPUT38), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n480), .A2(new_n486), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n493), .A2(new_n477), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n254), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n670), .A2(new_n448), .B1(G472), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n700), .B(new_n701), .C1(new_n672), .C2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n696), .A2(new_n698), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NAND2_X1  g522(.A1(new_n646), .A2(new_n680), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n636), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n673), .A2(new_n629), .A3(new_n684), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND4_X1  g526(.A1(new_n684), .A2(new_n264), .A3(new_n646), .A4(new_n629), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n586), .A2(new_n597), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n254), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n603), .A3(new_n254), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n561), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n513), .A2(new_n558), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT110), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n684), .A2(new_n264), .A3(new_n629), .A4(new_n656), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n720), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n280), .ZN(G18));
  NAND3_X1  g541(.A1(new_n513), .A2(new_n320), .A3(new_n665), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n684), .A2(new_n629), .A3(new_n719), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n357), .ZN(G21));
  NAND3_X1  g545(.A1(new_n684), .A2(new_n629), .A3(new_n699), .ZN(new_n732));
  OAI221_X1 g546(.A(new_n487), .B1(KEYINPUT31), .B2(new_n478), .C1(new_n477), .C2(new_n504), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n632), .A2(G472), .B1(new_n445), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n718), .A2(new_n263), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n558), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  AND3_X1   g552(.A1(new_n684), .A2(new_n629), .A3(new_n719), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n445), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n633), .A2(new_n665), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n709), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(G125), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G27));
  OAI211_X1 g559(.A(new_n439), .B(new_n443), .C1(new_n440), .C2(new_n441), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n607), .ZN(new_n747));
  INV_X1    g561(.A(new_n709), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n513), .A3(new_n558), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n557), .B1(new_n671), .B2(new_n672), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT42), .A3(new_n748), .A4(new_n747), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n751), .A2(KEYINPUT112), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n190), .ZN(G33));
  NOR2_X1   g573(.A1(new_n655), .A2(new_n681), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n747), .A2(new_n513), .A3(new_n558), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  INV_X1    g576(.A(new_n645), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n317), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(KEYINPUT114), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT114), .B(KEYINPUT43), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n766), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n635), .A2(new_n665), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT44), .Z(new_n770));
  OAI21_X1  g584(.A(new_n599), .B1(new_n601), .B2(new_n596), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT113), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n603), .B1(new_n771), .B2(new_n772), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n604), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n717), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n561), .B(new_n688), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n770), .A2(new_n746), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  INV_X1    g596(.A(new_n513), .ZN(new_n783));
  INV_X1    g597(.A(new_n746), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n558), .A2(new_n709), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n561), .B1(new_n778), .B2(new_n779), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(KEYINPUT47), .B(new_n561), .C1(new_n778), .C2(new_n779), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n201), .ZN(G42));
  INV_X1    g606(.A(new_n443), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n764), .A2(new_n560), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n716), .A2(new_n717), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n558), .B(new_n794), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT115), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n705), .A2(new_n672), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n797), .B2(new_n796), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n701), .A3(new_n801), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n729), .A2(new_n728), .B1(new_n732), .B2(new_n736), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n721), .A3(new_n726), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n253), .A2(new_n269), .A3(new_n307), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n645), .B1(new_n315), .B2(new_n316), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n805), .A2(new_n806), .A3(new_n264), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n442), .A2(new_n443), .A3(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n558), .A3(new_n661), .A4(new_n611), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n612), .A2(new_n666), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n651), .A2(new_n652), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n269), .A2(new_n811), .A3(new_n307), .A4(new_n680), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n608), .A2(new_n812), .A3(new_n610), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n746), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n513), .A3(new_n665), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n747), .A2(new_n665), .A3(new_n734), .A4(new_n748), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n761), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n804), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n758), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n626), .A2(new_n630), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n607), .A2(new_n681), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n669), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n705), .B2(new_n672), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n822), .A3(new_n699), .A4(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n665), .A2(new_n607), .A3(new_n681), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n512), .A2(KEYINPUT32), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n704), .A2(G472), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n500), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT116), .B1(new_n732), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n743), .A2(new_n685), .A3(new_n711), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT52), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n743), .A2(new_n685), .A3(new_n711), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n826), .A2(new_n832), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n819), .A2(new_n820), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n839), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n804), .A2(new_n756), .A3(new_n818), .A4(new_n757), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT117), .B1(new_n810), .B2(new_n817), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n841), .B1(new_n751), .B2(new_n753), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n804), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n817), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n612), .A2(new_n666), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n809), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n835), .A3(new_n839), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n845), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n847), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n674), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n768), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n768), .A2(KEYINPUT118), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n558), .A3(new_n734), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n701), .A2(new_n793), .A3(new_n719), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT50), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n867), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n746), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n789), .A2(new_n790), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n795), .A2(new_n561), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n864), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n784), .A2(new_n719), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n741), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n876), .A2(new_n800), .A3(new_n557), .A4(new_n262), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n763), .A2(new_n315), .A3(new_n316), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n877), .A2(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n870), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n879), .B2(new_n646), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT48), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n877), .B2(new_n752), .ZN(new_n889));
  INV_X1    g703(.A(new_n752), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n875), .A2(KEYINPUT48), .A3(new_n890), .A4(new_n876), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n865), .A2(KEYINPUT120), .A3(new_n729), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT120), .B1(new_n865), .B2(new_n729), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n858), .A2(new_n884), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n802), .B1(new_n897), .B2(new_n898), .ZN(G75));
  NAND2_X1  g713(.A1(new_n845), .A2(new_n856), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G902), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n369), .B(new_n416), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n255), .A2(G952), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT122), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n901), .A2(new_n440), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n905), .B2(KEYINPUT121), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(KEYINPUT121), .B2(new_n905), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n906), .A2(new_n912), .ZN(G51));
  INV_X1    g727(.A(new_n908), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n857), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n845), .A2(new_n856), .A3(KEYINPUT123), .A4(new_n848), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n604), .B(KEYINPUT57), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n714), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n902), .A2(new_n776), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n922), .B2(new_n923), .ZN(G54));
  NAND4_X1  g738(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n249), .A2(new_n250), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n908), .B1(new_n925), .B2(new_n928), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n925), .B2(new_n928), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G60));
  XNOR2_X1  g746(.A(new_n643), .B(KEYINPUT59), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n847), .B2(new_n857), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n639), .A2(new_n641), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n908), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n933), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n919), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(G63));
  XOR2_X1   g754(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n941));
  INV_X1    g755(.A(new_n843), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n804), .A2(new_n855), .A3(new_n849), .A4(new_n850), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n840), .A2(new_n841), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n549), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n663), .B(new_n946), .C1(new_n845), .C2(new_n856), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n947), .B(new_n908), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n946), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n900), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n952), .A2(KEYINPUT126), .A3(new_n663), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n941), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n908), .A3(new_n947), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n257), .B2(new_n411), .ZN(new_n959));
  NOR4_X1   g773(.A1(new_n810), .A2(new_n803), .A3(new_n721), .A4(new_n726), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n369), .B1(G898), .B2(new_n255), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n238), .A2(new_n239), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n484), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(G900), .A2(G953), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n780), .A2(new_n890), .A3(new_n732), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n791), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n761), .A3(new_n781), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n970), .A2(new_n758), .A3(new_n834), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n967), .B1(new_n971), .B2(new_n255), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n707), .A2(new_n836), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n707), .A2(new_n978), .A3(new_n836), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n805), .A2(new_n806), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n693), .A2(new_n752), .A3(new_n784), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n781), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n791), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n977), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n984), .A2(new_n255), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n973), .B(new_n975), .C1(new_n985), .C2(new_n965), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n965), .B1(new_n984), .B2(new_n255), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n974), .B1(new_n987), .B2(new_n972), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n842), .A2(new_n846), .ZN(new_n993));
  INV_X1    g807(.A(new_n702), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n502), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n971), .B2(new_n960), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n485), .B(KEYINPUT127), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(new_n477), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n908), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n477), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n977), .A2(new_n960), .A3(new_n979), .A4(new_n983), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n991), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n995), .A2(new_n999), .A3(new_n1002), .ZN(G57));
endmodule


