//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1336, new_n1337, new_n1338, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1410, new_n1411;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n202), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n209), .B(new_n213), .C1(G87), .C2(G250), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(G244), .Z(new_n215));
  AND2_X1   g0015(.A1(KEYINPUT64), .A2(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(KEYINPUT64), .A2(G68), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n215), .A2(G77), .B1(new_n218), .B2(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n214), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(G20), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n225), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G226), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n229), .ZN(new_n256));
  INV_X1    g0056(.A(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(G33), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n218), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n202), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n256), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT11), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT12), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n257), .A2(G1), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT72), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(new_n256), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n229), .A4(new_n255), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(G68), .B1(new_n275), .B2(new_n268), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT64), .A2(G68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT64), .A2(G68), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n279), .A2(KEYINPUT12), .A3(G20), .A4(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n265), .A2(new_n269), .A3(new_n276), .A4(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(KEYINPUT77), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  OAI211_X1 g0088(.A(G232), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT75), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT75), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(G232), .A4(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(G226), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G97), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n290), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G1), .A3(G13), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n302), .ZN(new_n305));
  INV_X1    g0105(.A(G238), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n286), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  AOI211_X1 g0109(.A(KEYINPUT13), .B(new_n307), .C1(new_n297), .C2(new_n300), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n285), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI221_X1 g0113(.A(G169), .B1(KEYINPUT77), .B2(new_n284), .C1(new_n309), .C2(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n301), .A2(new_n308), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT76), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n301), .A2(new_n286), .A3(new_n308), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n310), .B1(new_n309), .B2(KEYINPUT76), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n283), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT76), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT13), .ZN(new_n326));
  OAI21_X1  g0126(.A(G190), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n283), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n311), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n302), .A2(new_n303), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n299), .A2(new_n302), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n215), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G238), .A2(G1698), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n335), .B1(new_n221), .B2(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n287), .A2(new_n288), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n211), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n338), .A3(new_n300), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(G179), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n312), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(G20), .ZN(new_n345));
  OR2_X1    g0145(.A1(KEYINPUT15), .A2(G87), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT15), .A2(G87), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G20), .A2(G77), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n349), .C1(new_n350), .C2(new_n262), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n275), .A2(G77), .B1(new_n256), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT73), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n272), .A2(new_n258), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n270), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n255), .A2(new_n229), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT72), .B1(new_n357), .B2(new_n267), .ZN(new_n358));
  INV_X1    g0158(.A(new_n274), .ZN(new_n359));
  OAI211_X1 g0159(.A(G77), .B(new_n356), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n351), .A2(new_n256), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT73), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n341), .B(new_n343), .C1(new_n355), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n355), .A2(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n340), .A2(G200), .ZN(new_n366));
  INV_X1    g0166(.A(G190), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n340), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n331), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n291), .A2(G222), .A3(new_n294), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT69), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT69), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n291), .A2(new_n373), .A3(G222), .A4(new_n294), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n291), .A2(G223), .A3(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n291), .A2(new_n258), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n300), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n333), .A2(G226), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n304), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(G179), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT70), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT8), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(G58), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT71), .B(new_n384), .C1(new_n350), .C2(new_n382), .ZN(new_n385));
  OR4_X1    g0185(.A1(new_n382), .A2(new_n220), .A3(KEYINPUT71), .A4(KEYINPUT8), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n345), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n203), .A2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n261), .A2(G150), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n256), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n267), .A2(G50), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n256), .A2(new_n270), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n202), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n380), .A2(new_n312), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n381), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n380), .A2(G200), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n391), .A2(KEYINPUT9), .A3(new_n393), .A4(new_n397), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n378), .A2(G190), .A3(new_n379), .A4(new_n304), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI211_X1 g0205(.A(new_n392), .B(new_n396), .C1(new_n390), .C2(new_n256), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n406), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT74), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n398), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n402), .B(new_n405), .C1(new_n407), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n403), .A2(new_n404), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT74), .B1(new_n406), .B2(KEYINPUT9), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n398), .A2(new_n408), .A3(new_n409), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT10), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n402), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n401), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n272), .B1(new_n385), .B2(new_n386), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n385), .A2(new_n386), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n422), .B2(new_n395), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT7), .B1(new_n337), .B2(new_n257), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT3), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n344), .ZN(new_n426));
  NAND2_X1  g0226(.A1(KEYINPUT3), .A2(G33), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(KEYINPUT7), .A3(new_n257), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G159), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n262), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n277), .A2(G58), .A3(new_n278), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n226), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n434), .B2(G20), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(new_n435), .A3(KEYINPUT16), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(new_n256), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT16), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n201), .B1(new_n218), .B2(G58), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n439), .A2(new_n257), .B1(new_n431), .B2(new_n262), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n426), .A2(new_n257), .A3(new_n427), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT7), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n279), .B1(new_n443), .B2(new_n428), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n438), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n423), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  OR2_X1    g0247(.A1(G223), .A2(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n210), .A2(G1698), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n287), .C2(new_n288), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G87), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n332), .B1(new_n452), .B2(new_n300), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n299), .A2(G232), .A3(new_n302), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n312), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n299), .B1(new_n450), .B2(new_n451), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n457), .A2(new_n316), .A3(new_n454), .A4(new_n332), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n447), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(G179), .A3(new_n455), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n457), .A2(new_n332), .A3(new_n454), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(KEYINPUT78), .C1(new_n461), .C2(new_n312), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT18), .B1(new_n446), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(G190), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n461), .A2(new_n329), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n446), .A2(KEYINPUT17), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n445), .A2(new_n256), .A3(new_n436), .ZN(new_n468));
  INV_X1    g0268(.A(new_n420), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n421), .B2(new_n394), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n468), .A2(new_n466), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT17), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n470), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT18), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n459), .A4(new_n462), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n464), .A2(new_n467), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n370), .A2(new_n419), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  AND2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G264), .A3(new_n299), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G274), .A3(new_n482), .ZN(new_n488));
  INV_X1    g0288(.A(G250), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n426), .A2(new_n427), .B1(new_n489), .B2(new_n294), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n208), .A2(G1698), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(G33), .B2(G294), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n486), .B(new_n488), .C1(new_n492), .C2(new_n299), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT84), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI221_X1 g0295(.A(new_n491), .B1(G250), .B2(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G294), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n300), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(KEYINPUT84), .A3(new_n486), .A4(new_n488), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(new_n367), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n493), .A2(new_n329), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n257), .B(G87), .C1(new_n287), .C2(new_n288), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n291), .A2(new_n507), .A3(new_n257), .A4(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n345), .A2(G116), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n257), .A3(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT23), .B1(new_n211), .B2(G20), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AND4_X1   g0315(.A1(new_n504), .A2(new_n509), .A3(new_n510), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n506), .B2(new_n508), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n504), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n256), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n272), .A2(new_n256), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n344), .A2(G1), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n211), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n281), .A2(G20), .A3(new_n211), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT25), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n519), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n503), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n487), .A2(new_n482), .B1(new_n230), .B2(new_n298), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n498), .A2(new_n300), .B1(new_n531), .B2(G264), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT84), .B1(new_n532), .B2(new_n488), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n299), .B1(new_n496), .B2(new_n497), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n485), .A2(G264), .A3(new_n299), .ZN(new_n535));
  INV_X1    g0335(.A(new_n488), .ZN(new_n536));
  NOR4_X1   g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n494), .ZN(new_n537));
  OAI21_X1  g0337(.A(G169), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(G179), .A3(new_n488), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n529), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT85), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n529), .A3(KEYINPUT85), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n530), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n266), .A2(G45), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n299), .A2(G250), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n482), .A2(G274), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G116), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n287), .A2(new_n288), .B1(G244), .B2(new_n294), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G238), .A2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(new_n300), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n316), .ZN(new_n555));
  INV_X1    g0355(.A(new_n552), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n291), .B(new_n556), .C1(G244), .C2(new_n294), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n299), .B1(new_n557), .B2(new_n550), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n312), .B1(new_n558), .B2(new_n549), .ZN(new_n559));
  INV_X1    g0359(.A(G87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n207), .A3(new_n211), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n296), .A2(new_n257), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT19), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n257), .B(G68), .C1(new_n287), .C2(new_n288), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n259), .B2(new_n207), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n256), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n346), .A2(new_n347), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n520), .A2(new_n570), .A3(new_n522), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n272), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n567), .A2(new_n256), .B1(new_n272), .B2(new_n569), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT82), .B1(new_n576), .B2(new_n571), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n555), .B(new_n559), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n553), .A2(new_n300), .ZN(new_n579));
  INV_X1    g0379(.A(new_n549), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n329), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n520), .A2(G87), .A3(new_n522), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n568), .A2(new_n572), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n554), .A2(G190), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT21), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n589), .B(new_n521), .C1(new_n273), .C2(new_n274), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n272), .A2(new_n589), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n255), .A2(new_n229), .B1(G20), .B2(new_n589), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G283), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n257), .C1(G33), .C2(new_n207), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT20), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G303), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n426), .A2(new_n599), .A3(new_n427), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G257), .A2(G1698), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n212), .B2(G1698), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n300), .B(new_n600), .C1(new_n602), .C2(new_n337), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n485), .A2(G270), .A3(new_n299), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n488), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G169), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n588), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G116), .B(new_n522), .C1(new_n358), .C2(new_n359), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n592), .A2(new_n594), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n594), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n608), .A2(new_n613), .A3(new_n591), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(KEYINPUT21), .A3(G169), .A4(new_n605), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n603), .A2(new_n488), .A3(new_n604), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(G179), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n607), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n605), .A2(G200), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n598), .B(new_n620), .C1(new_n367), .C2(new_n605), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n621), .A2(new_n607), .A3(new_n615), .A4(new_n617), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n587), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n485), .A2(G257), .A3(new_n299), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n489), .B1(new_n426), .B2(new_n427), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  OAI21_X1  g0428(.A(G1698), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(G244), .B1(new_n287), .B2(new_n288), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n630), .A2(new_n628), .B1(G33), .B2(G283), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n294), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n626), .B1(new_n633), .B2(new_n300), .ZN(new_n634));
  AOI211_X1 g0434(.A(KEYINPUT79), .B(new_n329), .C1(new_n634), .C2(new_n488), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT79), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n628), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n632), .A2(new_n637), .A3(new_n593), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n291), .A2(G250), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n294), .B1(new_n639), .B2(KEYINPUT4), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n300), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n626), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n488), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n636), .B1(new_n643), .B2(G200), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n267), .A2(G97), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n523), .B2(new_n207), .ZN(new_n647));
  OAI21_X1  g0447(.A(G107), .B1(new_n424), .B2(new_n429), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT6), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n207), .A2(new_n211), .ZN(new_n650));
  NOR2_X1   g0450(.A1(G97), .A2(G107), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n211), .A2(KEYINPUT6), .A3(G97), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n261), .A2(G77), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n648), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n657), .B2(new_n256), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n641), .A2(G190), .A3(new_n488), .A4(new_n642), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n635), .A2(new_n644), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n443), .A2(new_n428), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(G107), .B1(G77), .B2(new_n261), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n357), .B1(new_n663), .B2(new_n655), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT80), .B1(new_n664), .B2(new_n647), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT80), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n643), .A2(G169), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n634), .A2(G179), .A3(new_n488), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n665), .A2(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT81), .B1(new_n661), .B2(new_n670), .ZN(new_n671));
  AOI211_X1 g0471(.A(new_n536), .B(new_n626), .C1(new_n633), .C2(new_n300), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT79), .B1(new_n672), .B2(new_n329), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n643), .A2(new_n636), .A3(G200), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n658), .A3(new_n659), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n657), .A2(new_n256), .ZN(new_n676));
  INV_X1    g0476(.A(new_n647), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n666), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AOI211_X1 g0478(.A(KEYINPUT80), .B(new_n647), .C1(new_n657), .C2(new_n256), .ZN(new_n679));
  AND4_X1   g0479(.A1(G179), .A2(new_n641), .A3(new_n488), .A4(new_n642), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n312), .B1(new_n634), .B2(new_n488), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n678), .A2(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT81), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n675), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n671), .A2(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n480), .A2(new_n545), .A3(new_n625), .A4(new_n685), .ZN(G372));
  NAND2_X1  g0486(.A1(new_n573), .A2(new_n574), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n576), .A2(KEYINPUT82), .A3(new_n571), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n559), .A2(new_n555), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n689), .A2(new_n690), .B1(new_n585), .B2(new_n584), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n658), .B1(new_n668), .B2(new_n669), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n578), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n670), .B2(new_n691), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n501), .A2(new_n502), .ZN(new_n698));
  INV_X1    g0498(.A(new_n529), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n587), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n541), .A2(new_n618), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n682), .A4(new_n675), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n480), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n367), .B1(new_n321), .B2(new_n322), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n311), .A2(new_n329), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n283), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n341), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n709));
  AND4_X1   g0509(.A1(new_n353), .A2(new_n360), .A3(new_n354), .A4(new_n361), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n342), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT86), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT86), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n365), .A2(new_n713), .A3(new_n342), .A4(new_n708), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n324), .B1(new_n707), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n471), .B(KEYINPUT17), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n460), .B1(new_n312), .B2(new_n461), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n474), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n475), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n474), .A2(new_n719), .A3(KEYINPUT18), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n412), .A2(new_n418), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n401), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n704), .A2(new_n726), .ZN(G369));
  NOR2_X1   g0527(.A1(new_n280), .A2(G20), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n266), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT27), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT27), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n731), .A3(new_n266), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(G213), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT87), .B(G343), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT88), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n545), .B1(new_n699), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n541), .ZN(new_n739));
  INV_X1    g0539(.A(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT89), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n737), .A2(new_n598), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n622), .B2(new_n624), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n607), .A2(new_n615), .A3(new_n617), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G330), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT89), .B(G330), .C1(new_n745), .C2(new_n747), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n742), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n618), .A2(new_n740), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n545), .A2(new_n755), .B1(new_n739), .B2(new_n737), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT90), .Z(G399));
  INV_X1    g0558(.A(new_n232), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G41), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n561), .A2(G116), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(G1), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n227), .B2(new_n761), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n703), .A2(new_n737), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(KEYINPUT29), .ZN(new_n767));
  INV_X1    g0567(.A(new_n530), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n675), .A2(new_n682), .A3(new_n586), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n540), .A2(new_n529), .A3(KEYINPUT85), .ZN(new_n770));
  AOI21_X1  g0570(.A(KEYINPUT85), .B1(new_n540), .B2(new_n529), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n768), .B(new_n769), .C1(new_n772), .C2(new_n746), .ZN(new_n773));
  INV_X1    g0573(.A(new_n692), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT26), .B1(new_n774), .B2(new_n587), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n670), .A2(new_n693), .A3(new_n691), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(new_n578), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n737), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n767), .B1(KEYINPUT29), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n532), .A2(new_n554), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n603), .A2(G179), .A3(new_n604), .A4(new_n488), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT91), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(new_n672), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n616), .A2(new_n532), .A3(new_n554), .A4(G179), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT91), .B1(new_n643), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT30), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n554), .B(KEYINPUT92), .Z(new_n790));
  AND3_X1   g0590(.A1(new_n493), .A2(new_n316), .A3(new_n605), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n790), .A2(new_n643), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT93), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n783), .A2(new_n672), .A3(KEYINPUT30), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT93), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(new_n796), .A3(new_n792), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT31), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n737), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n789), .A2(new_n795), .A3(new_n792), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n740), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n798), .A2(new_n800), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n685), .A2(new_n545), .A3(new_n625), .A4(new_n737), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G330), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n780), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n765), .B1(new_n808), .B2(G1), .ZN(G364));
  NAND2_X1  g0609(.A1(new_n728), .A2(G45), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n761), .A2(G1), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n748), .B2(new_n749), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n750), .A2(new_n813), .A3(new_n752), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n811), .B(KEYINPUT94), .Z(new_n815));
  AOI21_X1  g0615(.A(new_n229), .B1(G20), .B2(new_n312), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n257), .A2(G179), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n329), .A2(G190), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n211), .ZN(new_n821));
  NAND2_X1  g0621(.A1(G20), .A2(G179), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n822), .A2(new_n367), .A3(new_n329), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n367), .A2(new_n329), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n818), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n824), .A2(new_n202), .B1(new_n826), .B2(new_n560), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n822), .A2(new_n329), .A3(G190), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n821), .B(new_n827), .C1(G68), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G190), .A2(G200), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n818), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n831), .A2(KEYINPUT32), .A3(new_n431), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n367), .A2(G179), .A3(G200), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n257), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n832), .B1(G97), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT32), .B1(new_n831), .B2(new_n431), .ZN(new_n837));
  AND4_X1   g0637(.A1(new_n291), .A2(new_n829), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n822), .A2(new_n367), .A3(G200), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n822), .A2(G190), .A3(G200), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT95), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(KEYINPUT95), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT96), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(KEYINPUT96), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n838), .B1(new_n220), .B2(new_n840), .C1(new_n258), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n337), .B1(new_n834), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n831), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n851), .A2(G329), .B1(G326), .B2(new_n823), .ZN(new_n852));
  INV_X1    g0652(.A(new_n828), .ZN(new_n853));
  XOR2_X1   g0653(.A(KEYINPUT33), .B(G317), .Z(new_n854));
  OAI21_X1  g0654(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n850), .B(new_n855), .C1(G322), .C2(new_n839), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n826), .B(KEYINPUT97), .Z(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(G303), .B1(G311), .B2(new_n844), .ZN(new_n859));
  INV_X1    g0659(.A(G283), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n856), .B(new_n859), .C1(new_n860), .C2(new_n820), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n817), .B1(new_n848), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(G13), .A2(G33), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(G20), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n816), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n759), .A2(new_n291), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n228), .A2(new_n481), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n867), .B(new_n868), .C1(new_n253), .C2(new_n481), .ZN(new_n869));
  INV_X1    g0669(.A(G355), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n291), .A2(new_n232), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(G116), .B2(new_n232), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n862), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n748), .ZN(new_n874));
  INV_X1    g0674(.A(new_n865), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n814), .B1(new_n815), .B2(new_n876), .ZN(G396));
  AOI21_X1  g0677(.A(new_n737), .B1(new_n363), .B2(new_n355), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n712), .A2(new_n714), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n740), .A2(new_n365), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n364), .B2(new_n369), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n675), .A2(new_n682), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n746), .B1(new_n529), .B2(new_n540), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n691), .B1(new_n503), .B2(new_n529), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT26), .B1(new_n682), .B2(new_n587), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n578), .A3(new_n694), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n737), .B(new_n882), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT100), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT100), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n703), .A2(new_n891), .A3(new_n737), .A4(new_n882), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n879), .A2(new_n881), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n890), .A2(new_n892), .B1(new_n766), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(new_n806), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(new_n811), .ZN(new_n896));
  INV_X1    g0696(.A(new_n815), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n816), .A2(new_n863), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(G77), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT98), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(G137), .A2(new_n823), .B1(new_n839), .B2(G143), .ZN(new_n903));
  INV_X1    g0703(.A(G150), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n903), .B1(new_n904), .B2(new_n853), .C1(new_n847), .C2(new_n431), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT34), .ZN(new_n906));
  INV_X1    g0706(.A(G132), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n291), .B1(new_n831), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n858), .B2(G50), .ZN(new_n909));
  INV_X1    g0709(.A(G68), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n820), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(G58), .B2(new_n835), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n337), .B1(new_n857), .B2(new_n211), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT99), .Z(new_n915));
  INV_X1    g0715(.A(new_n847), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(G116), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n835), .A2(G97), .B1(G311), .B2(new_n851), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n820), .A2(new_n560), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n824), .A2(new_n599), .B1(new_n840), .B2(new_n849), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(G283), .C2(new_n828), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n915), .A2(new_n917), .A3(new_n918), .A4(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n817), .B1(new_n913), .B2(new_n922), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n902), .B(new_n923), .C1(new_n863), .C2(new_n893), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n896), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(G384));
  NOR2_X1   g0726(.A1(KEYINPUT103), .A2(KEYINPUT31), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n802), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n801), .A2(new_n740), .A3(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n804), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(G179), .B1(new_n325), .B2(new_n326), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n313), .A3(new_n314), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n283), .B(new_n740), .C1(new_n707), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n740), .A2(new_n283), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n324), .A2(new_n330), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n893), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT101), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n910), .B1(new_n443), .B2(new_n428), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n438), .B1(new_n440), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n256), .A3(new_n436), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n470), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n939), .B1(new_n943), .B2(new_n734), .ZN(new_n944));
  AOI211_X1 g0744(.A(KEYINPUT101), .B(new_n733), .C1(new_n942), .C2(new_n470), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n477), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n474), .A2(new_n734), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT37), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n948), .A2(new_n949), .A3(new_n471), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n474), .A2(new_n459), .A3(new_n462), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n944), .A2(new_n945), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n943), .A2(new_n719), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n955), .A2(new_n471), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n949), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n947), .B(KEYINPUT38), .C1(new_n953), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n471), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n960), .A2(new_n945), .A3(new_n944), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n952), .B1(new_n961), .B2(new_n949), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n962), .B2(new_n947), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n932), .B(new_n938), .C1(new_n959), .C2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT38), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n948), .B1(new_n717), .B2(new_n723), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n720), .A2(new_n948), .A3(new_n471), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n950), .A2(new_n951), .B1(new_n969), .B2(KEYINPUT37), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n958), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n972), .A2(new_n932), .A3(KEYINPUT40), .A4(new_n938), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT104), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT40), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n958), .B2(new_n971), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT104), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(new_n977), .A3(new_n932), .A4(new_n938), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n966), .A2(new_n974), .A3(G330), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n480), .A2(G330), .A3(new_n932), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT105), .Z(new_n982));
  AND2_X1   g0782(.A1(new_n974), .A2(new_n978), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n983), .A2(new_n480), .A3(new_n932), .A4(new_n966), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n711), .A2(new_n740), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n890), .B2(new_n892), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n935), .A2(new_n937), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n959), .C2(new_n963), .ZN(new_n990));
  INV_X1    g0790(.A(new_n963), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(KEYINPUT39), .A3(new_n958), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT39), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n972), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n934), .A2(new_n283), .A3(new_n737), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n721), .A2(new_n722), .A3(new_n733), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n990), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n779), .A2(KEYINPUT29), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n480), .B1(new_n1000), .B2(new_n767), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n726), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n999), .B(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n985), .B(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n266), .B2(new_n728), .ZN(new_n1005));
  OAI211_X1 g0805(.A(G20), .B(new_n230), .C1(new_n654), .C2(KEYINPUT35), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n589), .B(new_n1006), .C1(KEYINPUT35), .C2(new_n654), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT36), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n228), .A2(G77), .A3(new_n433), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(G50), .B2(new_n910), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(G1), .A3(new_n280), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(new_n1008), .A3(new_n1011), .ZN(G367));
  XNOR2_X1  g0812(.A(new_n760), .B(KEYINPUT41), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n750), .A2(KEYINPUT110), .A3(new_n752), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n545), .A2(new_n755), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n742), .C2(new_n755), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n742), .B2(new_n755), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1017), .A2(KEYINPUT110), .A3(new_n750), .A4(new_n752), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1016), .A2(new_n780), .A3(new_n1018), .A4(new_n806), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n692), .A2(new_n740), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n737), .A2(new_n658), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n883), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT109), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n756), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT109), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1023), .B(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1028), .A2(KEYINPUT45), .A3(new_n756), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT44), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1028), .B2(new_n756), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1024), .A2(new_n1025), .A3(KEYINPUT44), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT111), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n754), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n754), .A2(new_n1036), .ZN(new_n1038));
  OAI211_X1 g0838(.A(KEYINPUT111), .B(new_n742), .C1(new_n751), .C2(new_n753), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n1034), .A4(new_n1030), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1019), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1013), .B1(new_n1041), .B2(new_n807), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n810), .A2(G1), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1015), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1028), .A2(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1047), .A2(KEYINPUT42), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(KEYINPUT42), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n670), .B1(new_n1028), .B2(new_n772), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1048), .B(new_n1049), .C1(new_n740), .C2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n737), .B1(new_n576), .B2(new_n582), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(new_n587), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT106), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n689), .A3(new_n690), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(KEYINPUT106), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT43), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1051), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n754), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT107), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1028), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1066), .B1(new_n1060), .B2(new_n1028), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1059), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n754), .A2(new_n1024), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1066), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1073), .A2(new_n1058), .A3(new_n1051), .A4(new_n1067), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1045), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n820), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(G97), .B1(new_n828), .B2(G294), .ZN(new_n1079));
  INV_X1    g0879(.A(G311), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1079), .B1(new_n599), .B2(new_n840), .C1(new_n1080), .C2(new_n824), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n291), .B(new_n1081), .C1(G107), .C2(new_n835), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n916), .A2(G283), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G317), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT46), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n858), .B2(G116), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n826), .A2(KEYINPUT46), .A3(new_n589), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1084), .B1(new_n1085), .B2(new_n831), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n826), .A2(new_n220), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n916), .A2(G50), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n834), .A2(new_n910), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G143), .B2(new_n823), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n904), .B2(new_n840), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT112), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  INV_X1    g0897(.A(G137), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n853), .A2(new_n431), .B1(new_n831), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n337), .B(new_n1099), .C1(G77), .C2(new_n1078), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1091), .A2(new_n1096), .A3(new_n1097), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1089), .B1(new_n1090), .B2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT47), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n815), .B1(new_n1103), .B2(new_n816), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n867), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n866), .B1(new_n232), .B2(new_n569), .C1(new_n244), .C2(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1057), .A2(new_n875), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1077), .A2(new_n1108), .ZN(G387));
  NAND2_X1  g0909(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n807), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n760), .A3(new_n1019), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1078), .A2(G116), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n291), .B1(new_n851), .B2(G326), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G322), .A2(new_n823), .B1(new_n828), .B2(G311), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n1085), .B2(new_n840), .C1(new_n847), .C2(new_n599), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT48), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n860), .B2(new_n834), .C1(new_n849), .C2(new_n826), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT49), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(KEYINPUT49), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1113), .B(new_n1114), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n834), .A2(new_n569), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n826), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G77), .A2(new_n1123), .B1(new_n851), .B2(G150), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n202), .B2(new_n840), .C1(new_n431), .C2(new_n824), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1122), .B(new_n1125), .C1(G68), .C2(new_n844), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1078), .A2(G97), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n422), .A2(new_n828), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1126), .A2(new_n291), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(KEYINPUT113), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT113), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n817), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n866), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n867), .B1(new_n241), .B2(new_n481), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n762), .B2(new_n871), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n350), .A2(G50), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G116), .B(new_n561), .C1(new_n1138), .C2(KEYINPUT50), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(G68), .A2(G77), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1138), .A2(KEYINPUT50), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1139), .A2(new_n481), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1137), .A2(new_n1142), .B1(new_n211), .B2(new_n759), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n897), .B1(new_n1135), .B2(new_n1143), .C1(new_n742), .C2(new_n875), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1112), .B1(new_n1044), .B2(new_n1110), .C1(new_n1134), .C2(new_n1144), .ZN(G393));
  NAND2_X1  g0945(.A1(new_n851), .A2(G143), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n202), .B2(new_n853), .C1(new_n279), .C2(new_n826), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n337), .B(new_n1147), .C1(G77), .C2(new_n835), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n824), .A2(new_n904), .B1(new_n840), .B2(new_n431), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT51), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n919), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1148), .B(new_n1153), .C1(new_n350), .C2(new_n847), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT114), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n851), .A2(G322), .B1(G303), .B2(new_n828), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n211), .B2(new_n820), .C1(new_n860), .C2(new_n826), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n291), .B(new_n1157), .C1(G116), .C2(new_n835), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n844), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n849), .B2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G317), .A2(new_n823), .B1(new_n839), .B2(G311), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT52), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1155), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT115), .Z(new_n1164));
  AOI21_X1  g0964(.A(new_n815), .B1(new_n1164), .B2(new_n816), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n248), .A2(new_n867), .B1(G97), .B2(new_n759), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n866), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1024), .A2(new_n865), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(new_n1043), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1037), .A2(new_n1040), .A3(new_n1019), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n760), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1173), .B2(new_n1041), .ZN(G390));
  INV_X1    g0974(.A(new_n989), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n995), .B1(new_n987), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n992), .A2(new_n994), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n778), .A2(new_n737), .A3(new_n882), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n986), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n989), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n996), .B1(new_n958), .B2(new_n971), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n932), .A2(new_n938), .A3(G330), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n893), .A2(new_n749), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n803), .B2(new_n804), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n989), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1178), .A2(new_n1184), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n989), .B1(new_n932), .B2(new_n1188), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1181), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1186), .B1(new_n1190), .B2(new_n989), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n988), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT116), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT116), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n988), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1194), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n980), .B(new_n726), .C1(new_n780), .C2(new_n479), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1187), .B(new_n1192), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1201), .ZN(new_n1203));
  OR3_X1    g1003(.A1(new_n1191), .A2(new_n1181), .A3(new_n1193), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1195), .A2(new_n988), .A3(new_n1198), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1198), .B1(new_n1195), .B2(new_n988), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1178), .A2(new_n1184), .A3(new_n1191), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1186), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1203), .B(new_n1207), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1202), .A2(new_n1211), .A3(new_n760), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1177), .A2(new_n863), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n421), .A2(new_n898), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n916), .A2(G97), .B1(G107), .B2(new_n828), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n860), .B2(new_n824), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT117), .Z(new_n1217));
  OAI21_X1  g1017(.A(new_n337), .B1(new_n857), .B2(new_n560), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT118), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n911), .B(new_n1219), .C1(G116), .C2(new_n839), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n835), .A2(G77), .B1(G294), .B2(new_n851), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1217), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n840), .A2(new_n907), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1078), .A2(G50), .B1(new_n828), .B2(G137), .ZN(new_n1224));
  INV_X1    g1024(.A(G125), .ZN(new_n1225));
  INV_X1    g1025(.A(G128), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n831), .C1(new_n1226), .C2(new_n824), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n337), .B(new_n1227), .C1(G159), .C2(new_n835), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT54), .B(G143), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n916), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n826), .A2(new_n904), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT53), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1222), .B1(new_n1223), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n815), .B1(new_n1234), .B2(new_n816), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1213), .A2(new_n1214), .A3(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT119), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1176), .A2(new_n1177), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1192), .B1(new_n1238), .B2(new_n1209), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1043), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1212), .A2(new_n1240), .ZN(G378));
  INV_X1    g1041(.A(G41), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G50), .B1(new_n427), .B2(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G58), .A2(new_n1078), .B1(new_n851), .B2(G283), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n258), .B2(new_n826), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1245), .A2(G41), .A3(new_n291), .A4(new_n1092), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n824), .A2(new_n589), .B1(new_n840), .B2(new_n211), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n570), .B2(new_n844), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(new_n207), .C2(new_n853), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1249), .B(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n824), .A2(new_n1225), .B1(new_n853), .B2(new_n907), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1123), .B2(new_n1229), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n904), .B2(new_n834), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G137), .B2(new_n844), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1226), .B2(new_n840), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT59), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G33), .B1(new_n1078), .B2(G159), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G41), .B1(new_n851), .B2(G124), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1243), .B(new_n1252), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n812), .B1(new_n1263), .B2(new_n817), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT122), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT55), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n419), .A2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(KEYINPUT55), .B(new_n401), .C1(new_n412), .C2(new_n418), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n398), .A2(new_n734), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n417), .B1(new_n416), .B2(new_n402), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n400), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT55), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n419), .A2(new_n1266), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1265), .B1(new_n1272), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1271), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1278), .A3(new_n1273), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(KEYINPUT122), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1264), .B1(new_n1284), .B2(new_n863), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n898), .A2(new_n202), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n983), .A2(new_n1284), .A3(G330), .A4(new_n966), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n990), .A2(new_n997), .A3(new_n998), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1272), .A2(new_n1279), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n979), .A2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1294), .B2(new_n1044), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n979), .A2(new_n1290), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1281), .A2(new_n1282), .A3(KEYINPUT122), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT122), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n979), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n999), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1211), .A2(new_n1203), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n761), .B1(new_n1303), .B2(KEYINPUT57), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT57), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1201), .B1(new_n1239), .B2(new_n1207), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1294), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1295), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(G375));
  NAND2_X1  g1109(.A1(new_n1207), .A2(new_n1203), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1204), .B(new_n1201), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1013), .A3(new_n1311), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1229), .A2(new_n828), .B1(new_n823), .B2(G132), .ZN(new_n1313));
  OAI221_X1 g1113(.A(new_n1313), .B1(new_n1226), .B2(new_n831), .C1(new_n1098), .C2(new_n840), .ZN(new_n1314));
  AOI211_X1 g1114(.A(new_n337), .B(new_n1314), .C1(G50), .C2(new_n835), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n858), .A2(G159), .B1(G150), .B2(new_n844), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1315), .B(new_n1316), .C1(new_n220), .C2(new_n820), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(G116), .A2(new_n828), .B1(new_n839), .B2(G283), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n599), .B2(new_n831), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1122), .B(new_n1319), .C1(G294), .C2(new_n823), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n1320), .B1(new_n207), .B2(new_n857), .C1(new_n211), .C2(new_n847), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n337), .B1(new_n820), .B2(new_n258), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(KEYINPUT123), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1317), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n815), .B1(new_n1324), .B2(new_n816), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n989), .B2(new_n864), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n910), .B2(new_n898), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1207), .B2(new_n1043), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1312), .A2(new_n1328), .ZN(G381));
  XNOR2_X1  g1129(.A(new_n1308), .B(KEYINPUT124), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(G378), .ZN(new_n1331));
  INV_X1    g1131(.A(G390), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1077), .A2(new_n1108), .A3(new_n1332), .ZN(new_n1333));
  NOR4_X1   g1133(.A1(new_n1333), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1331), .A2(new_n925), .A3(new_n1334), .ZN(G407));
  INV_X1    g1135(.A(G213), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n735), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1331), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(G407), .ZN(G409));
  NAND2_X1  g1139(.A1(new_n1211), .A2(new_n1203), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(KEYINPUT57), .A3(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1307), .A2(new_n1342), .A3(new_n760), .ZN(new_n1343));
  AOI22_X1  g1143(.A1(new_n1341), .A2(new_n1043), .B1(new_n1286), .B2(new_n1285), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(G378), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1303), .A2(new_n1013), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1344), .ZN(new_n1347));
  INV_X1    g1147(.A(G378), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1345), .A2(new_n1349), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n735), .A2(new_n1336), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT125), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT60), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1311), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1356), .A2(KEYINPUT60), .A3(new_n1201), .A4(new_n1204), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1355), .A2(new_n1357), .A3(new_n1310), .A4(new_n760), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1328), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1353), .B1(new_n1359), .B2(new_n925), .ZN(new_n1360));
  AOI211_X1 g1160(.A(KEYINPUT125), .B(G384), .C1(new_n1358), .C2(new_n1328), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1358), .A2(G384), .A3(new_n1328), .ZN(new_n1362));
  NOR3_X1   g1162(.A1(new_n1360), .A2(new_n1361), .A3(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1350), .A2(new_n1352), .A3(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1364), .A2(KEYINPUT62), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1351), .A2(G2897), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1362), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1367), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1370));
  NOR4_X1   g1170(.A1(new_n1360), .A2(new_n1361), .A3(new_n1366), .A4(new_n1362), .ZN(new_n1371));
  AOI21_X1  g1171(.A(G378), .B1(new_n1346), .B2(new_n1344), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1372), .B1(new_n1308), .B2(G378), .ZN(new_n1373));
  OAI22_X1  g1173(.A1(new_n1370), .A2(new_n1371), .B1(new_n1373), .B2(new_n1351), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT61), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT62), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1350), .A2(new_n1376), .A3(new_n1352), .A4(new_n1363), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1365), .A2(new_n1374), .A3(new_n1375), .A4(new_n1377), .ZN(new_n1378));
  XOR2_X1   g1178(.A(G393), .B(G396), .Z(new_n1379));
  AOI21_X1  g1179(.A(new_n1332), .B1(new_n1077), .B2(new_n1108), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1075), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1108), .ZN(new_n1382));
  NOR3_X1   g1182(.A1(new_n1381), .A2(new_n1382), .A3(G390), .ZN(new_n1383));
  OAI21_X1  g1183(.A(new_n1379), .B1(new_n1380), .B2(new_n1383), .ZN(new_n1384));
  OAI21_X1  g1184(.A(G390), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1385));
  XNOR2_X1  g1185(.A(G393), .B(G396), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1333), .A2(new_n1385), .A3(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1384), .A2(new_n1387), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1378), .A2(new_n1388), .ZN(new_n1389));
  INV_X1    g1189(.A(KEYINPUT126), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1364), .A2(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1391), .A2(KEYINPUT63), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1363), .A2(new_n1367), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1359), .A2(new_n925), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1394), .A2(KEYINPUT125), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1359), .A2(new_n925), .A3(new_n1353), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1395), .A2(new_n1369), .A3(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1397), .A2(new_n1366), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1393), .A2(new_n1398), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(new_n1350), .A2(new_n1352), .ZN(new_n1400));
  NAND3_X1  g1200(.A1(new_n1384), .A2(new_n1375), .A3(new_n1387), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1401), .A2(KEYINPUT127), .ZN(new_n1402));
  INV_X1    g1202(.A(KEYINPUT127), .ZN(new_n1403));
  NAND4_X1  g1203(.A1(new_n1384), .A2(new_n1403), .A3(new_n1375), .A4(new_n1387), .ZN(new_n1404));
  AOI22_X1  g1204(.A1(new_n1399), .A2(new_n1400), .B1(new_n1402), .B2(new_n1404), .ZN(new_n1405));
  INV_X1    g1205(.A(KEYINPUT63), .ZN(new_n1406));
  NAND3_X1  g1206(.A1(new_n1364), .A2(new_n1390), .A3(new_n1406), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1392), .A2(new_n1405), .A3(new_n1407), .ZN(new_n1408));
  NAND2_X1  g1208(.A1(new_n1389), .A2(new_n1408), .ZN(G405));
  XNOR2_X1  g1209(.A(new_n1388), .B(new_n1363), .ZN(new_n1410));
  XNOR2_X1  g1210(.A(new_n1308), .B(G378), .ZN(new_n1411));
  XNOR2_X1  g1211(.A(new_n1410), .B(new_n1411), .ZN(G402));
endmodule


