//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972;
  NOR2_X1   g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT94), .B(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G43gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(KEYINPUT95), .A3(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT95), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n216));
  MUX2_X1   g015(.A(new_n207), .B(new_n215), .S(new_n216), .Z(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT17), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(G8gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT96), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(new_n223), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n217), .B(new_n223), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n228), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n228), .A3(new_n226), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G197gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT11), .B(G169gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n229), .A2(new_n243), .A3(new_n232), .A4(new_n235), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G141gat), .B(G148gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(G155gat), .B2(G162gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G141gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G148gat), .ZN(new_n255));
  INV_X1    g054(.A(G148gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G141gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G155gat), .B(G162gat), .ZN(new_n259));
  INV_X1    g058(.A(G155gat), .ZN(new_n260));
  INV_X1    g059(.A(G162gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT2), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n253), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n253), .A2(new_n263), .A3(KEYINPUT76), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G197gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G197gat), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n276), .A2(new_n278), .A3(G204gat), .ZN(new_n279));
  AOI21_X1  g078(.A(G204gat), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(G211gat), .A2(G218gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n283));
  NAND2_X1  g082(.A1(G211gat), .A2(G218gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n274), .C1(new_n279), .C2(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n271), .A2(new_n272), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G228gat), .A2(G233gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n267), .B2(new_n268), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT83), .B1(new_n294), .B2(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n253), .A2(new_n263), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G204gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n277), .A2(G197gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n276), .A2(new_n278), .A3(G204gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n273), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(new_n285), .ZN(new_n305));
  INV_X1    g104(.A(new_n288), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n270), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT3), .B1(new_n307), .B2(KEYINPUT82), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT29), .B1(new_n287), .B2(new_n288), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n298), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n282), .A2(new_n284), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n281), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316));
  INV_X1    g115(.A(new_n314), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n274), .C1(new_n279), .C2(new_n280), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n315), .A2(new_n316), .A3(new_n270), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n264), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n281), .B2(new_n314), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n316), .B1(new_n321), .B2(new_n318), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n297), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n289), .B1(new_n269), .B2(new_n270), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n293), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT84), .B1(new_n313), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n325), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n292), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n264), .B1(new_n309), .B2(new_n310), .ZN(new_n330));
  AOI211_X1 g129(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n287), .C2(new_n288), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n297), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n293), .A3(new_n291), .A4(new_n295), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(G22gat), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n327), .A2(new_n335), .A3(KEYINPUT85), .A4(G22gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G78gat), .B(G106gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(G50gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n270), .B1(new_n304), .B2(new_n317), .ZN(new_n345));
  INV_X1    g144(.A(new_n318), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT81), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n264), .A3(new_n319), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n324), .B1(new_n348), .B2(new_n297), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n296), .A2(new_n312), .B1(new_n349), .B2(new_n293), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n344), .B1(new_n350), .B2(G22gat), .ZN(new_n351));
  INV_X1    g150(.A(G22gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n329), .A2(new_n333), .A3(KEYINPUT86), .A4(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n343), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n350), .A2(G22gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n329), .B2(new_n333), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n343), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n355), .A2(KEYINPUT87), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT87), .B1(new_n355), .B2(new_n358), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT69), .B(G113gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G120gat), .ZN(new_n362));
  INV_X1    g161(.A(G134gat), .ZN(new_n363));
  INV_X1    g162(.A(G127gat), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT70), .B(G127gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G134gat), .ZN(new_n369));
  INV_X1    g168(.A(G113gat), .ZN(new_n370));
  INV_X1    g169(.A(G120gat), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT1), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n362), .A2(new_n367), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(KEYINPUT67), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G134gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n376), .A3(G127gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT68), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G127gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n381), .B2(new_n363), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n372), .B1(new_n370), .B2(new_n371), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT4), .B1(new_n385), .B2(new_n297), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n298), .A2(new_n387), .A3(new_n373), .A4(new_n384), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(KEYINPUT79), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n269), .B(new_n385), .C1(new_n264), .C2(new_n298), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n391), .B(KEYINPUT4), .C1(new_n385), .C2(new_n297), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n385), .B(new_n298), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n394), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n386), .A2(new_n388), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(new_n401), .A3(new_n394), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n385), .B(new_n297), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT77), .A3(new_n395), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n400), .A2(new_n402), .A3(new_n404), .A4(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n405), .A3(new_n411), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n412), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT23), .ZN(new_n420));
  NAND2_X1  g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(G169gat), .B2(G176gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT64), .ZN(new_n426));
  INV_X1    g225(.A(G183gat), .ZN(new_n427));
  INV_X1    g226(.A(G190gat), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT24), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT24), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(G183gat), .A3(G190gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n424), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n425), .B1(new_n429), .B2(new_n431), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n420), .A2(KEYINPUT25), .A3(new_n423), .A4(new_n421), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n433), .A2(KEYINPUT25), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT27), .B(G183gat), .Z(new_n437));
  OAI21_X1  g236(.A(KEYINPUT28), .B1(new_n437), .B2(G190gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT66), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT65), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n439), .B(G183gat), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT65), .B(KEYINPUT27), .C1(new_n427), .C2(KEYINPUT66), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n441), .B2(G183gat), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(G169gat), .B2(G176gat), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n419), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n438), .A2(new_n446), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n436), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G226gat), .A2(G233gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n452), .B(KEYINPUT75), .Z(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n436), .B2(new_n450), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n290), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n434), .A2(new_n435), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n426), .A2(new_n432), .ZN(new_n458));
  INV_X1    g257(.A(new_n424), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT25), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n450), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n453), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n452), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n464), .B(new_n289), .C1(new_n465), .C2(new_n451), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n456), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G8gat), .B(G36gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  OR3_X1    g270(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n270), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  INV_X1    g272(.A(new_n453), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n455), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n289), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n466), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n456), .A2(new_n466), .A3(new_n470), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n418), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n359), .A2(new_n360), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  INV_X1    g285(.A(new_n385), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n462), .B2(new_n463), .ZN(new_n488));
  INV_X1    g287(.A(G227gat), .ZN(new_n489));
  INV_X1    g288(.A(G233gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n436), .A2(new_n385), .A3(new_n450), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT32), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT33), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G15gat), .B(G43gat), .Z(new_n497));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n499), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n493), .B(KEYINPUT32), .C1(new_n495), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n492), .ZN(new_n505));
  INV_X1    g304(.A(new_n491), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g306(.A(KEYINPUT34), .B(new_n491), .C1(new_n488), .C2(new_n492), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n500), .A3(new_n502), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT71), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n500), .A3(new_n502), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT72), .B(new_n486), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n509), .A2(new_n500), .A3(new_n502), .ZN(new_n518));
  INV_X1    g317(.A(new_n507), .ZN(new_n519));
  INV_X1    g318(.A(new_n508), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n500), .A2(new_n502), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n518), .B2(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n515), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT72), .B1(new_n527), .B2(new_n486), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT88), .B1(new_n485), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n355), .A2(new_n358), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n418), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n482), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n355), .A2(KEYINPUT87), .A3(new_n358), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n486), .B1(new_n513), .B2(new_n516), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(new_n523), .A3(new_n517), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT89), .B(KEYINPUT39), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n393), .A2(new_n395), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n411), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT39), .B1(new_n403), .B2(new_n395), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n393), .B2(new_n395), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n393), .A2(new_n395), .ZN(new_n552));
  INV_X1    g351(.A(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(KEYINPUT90), .A3(new_n411), .A4(new_n546), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n550), .A2(new_n555), .A3(KEYINPUT91), .A4(new_n551), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n554), .A2(KEYINPUT40), .A3(new_n411), .A4(new_n546), .ZN(new_n561));
  AND4_X1   g360(.A1(new_n413), .A2(new_n472), .A3(new_n481), .A4(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n476), .B(new_n289), .C1(new_n453), .C2(new_n451), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n564), .A2(KEYINPUT92), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n464), .B1(new_n451), .B2(new_n465), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n564), .A2(KEYINPUT92), .B1(new_n566), .B2(new_n290), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT38), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n569), .B(new_n471), .C1(new_n467), .C2(KEYINPUT37), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n480), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n471), .A2(KEYINPUT37), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n479), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n467), .A2(KEYINPUT37), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n560), .A2(new_n562), .B1(new_n418), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n359), .B2(new_n360), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n530), .A2(new_n543), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n359), .A2(new_n360), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n535), .A2(new_n527), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n484), .B(new_n522), .C1(new_n359), .C2(new_n360), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n246), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G57gat), .A2(G64gat), .ZN(new_n589));
  OR2_X1    g388(.A1(G57gat), .A2(G64gat), .ZN(new_n590));
  INV_X1    g389(.A(G71gat), .ZN(new_n591));
  INV_X1    g390(.A(G78gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n589), .B(new_n590), .C1(new_n593), .C2(KEYINPUT9), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT97), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n592), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n594), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT20), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n223), .B1(KEYINPUT21), .B2(new_n599), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT99), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G99gat), .B(G106gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n218), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n217), .A2(new_n623), .B1(KEYINPUT41), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT101), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n628), .B(new_n630), .Z(new_n631));
  NOR2_X1   g430(.A1(new_n626), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT100), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n628), .B(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n614), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n623), .B(new_n598), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(KEYINPUT102), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n599), .A2(new_n623), .A3(KEYINPUT10), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT102), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n644), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n653), .A2(KEYINPUT103), .A3(new_n646), .A4(new_n645), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n643), .A2(new_n650), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n646), .A3(new_n645), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n650), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n656), .ZN(new_n663));
  INV_X1    g462(.A(new_n659), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT104), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n641), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n588), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n534), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(G1gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  OAI21_X1  g476(.A(G8gat), .B1(new_n673), .B2(new_n482), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT106), .B(KEYINPUT16), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G8gat), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n588), .A2(new_n483), .A3(new_n672), .A4(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n677), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT107), .ZN(G1325gat));
  OAI21_X1  g483(.A(KEYINPUT108), .B1(new_n524), .B2(new_n528), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n541), .A2(new_n686), .A3(new_n523), .A4(new_n517), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n673), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n527), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n673), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n588), .A2(new_n580), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n671), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(new_n640), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n579), .B2(new_n587), .ZN(new_n697));
  INV_X1    g496(.A(new_n670), .ZN(new_n698));
  INV_X1    g497(.A(new_n614), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n246), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n206), .A3(new_n418), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n579), .A2(new_n587), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n640), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n537), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n533), .A2(KEYINPUT109), .A3(new_n535), .A4(new_n536), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n688), .A2(new_n713), .A3(new_n578), .A4(new_n714), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n696), .B(new_n711), .C1(new_n715), .C2(new_n587), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n702), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n534), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n706), .A2(new_n719), .ZN(G1328gat));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n205), .A3(new_n483), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  NOR2_X1   g521(.A1(new_n718), .A2(new_n482), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n205), .B2(new_n723), .ZN(G1329gat));
  NOR3_X1   g523(.A1(new_n703), .A2(G43gat), .A3(new_n527), .ZN(new_n725));
  INV_X1    g524(.A(new_n688), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n717), .A2(new_n726), .A3(new_n702), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(G43gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT47), .ZN(G1330gat));
  NOR4_X1   g528(.A1(new_n692), .A2(G50gat), .A3(new_n696), .A4(new_n701), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n717), .A2(new_n580), .A3(new_n702), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(G50gat), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT111), .B1(new_n731), .B2(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI221_X4 g534(.A(new_n730), .B1(KEYINPUT111), .B2(KEYINPUT48), .C1(new_n731), .C2(G50gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  NAND2_X1  g536(.A1(new_n715), .A2(new_n587), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n246), .A2(new_n738), .A3(new_n641), .A4(new_n698), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n418), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n483), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(new_n527), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n739), .A2(new_n591), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n739), .A2(new_n726), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n591), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n580), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g551(.A1(new_n699), .A2(new_n245), .A3(new_n670), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n717), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n618), .B1(new_n754), .B2(new_n418), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n699), .A2(new_n245), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n714), .A2(new_n578), .A3(new_n685), .A4(new_n687), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n485), .A2(KEYINPUT109), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n581), .A2(new_n583), .B1(new_n585), .B2(KEYINPUT35), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n640), .B(new_n756), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n640), .A4(new_n756), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n698), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(G85gat), .A3(new_n534), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n755), .A2(new_n767), .ZN(G1336gat));
  NOR2_X1   g567(.A1(new_n482), .A2(G92gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n670), .B(new_n770), .C1(new_n763), .C2(new_n764), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n483), .B(new_n753), .C1(new_n709), .C2(new_n716), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n771), .B1(new_n775), .B2(KEYINPUT112), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n778), .A3(G92gat), .ZN(new_n779));
  AOI211_X1 g578(.A(KEYINPUT113), .B(new_n773), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n775), .A2(KEYINPUT112), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n779), .A3(new_n772), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n781), .B1(new_n783), .B2(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n776), .B1(new_n780), .B2(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n754), .B2(new_n726), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n766), .A2(G99gat), .A3(new_n527), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(new_n788), .ZN(G1338gat));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n754), .A2(new_n580), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n581), .A2(G106gat), .A3(new_n670), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT114), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n791), .A2(G106gat), .B1(new_n765), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n791), .A2(G106gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n790), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n790), .A2(new_n794), .B1(new_n795), .B2(new_n797), .ZN(G1339gat));
  NOR2_X1   g597(.A1(new_n671), .A2(new_n245), .ZN(new_n799));
  INV_X1    g598(.A(new_n650), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n653), .A2(new_n800), .A3(new_n646), .A4(new_n645), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n655), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n661), .A2(new_n803), .A3(new_n650), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n664), .A4(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n800), .B1(new_n661), .B2(new_n642), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n654), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n664), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(new_n811), .A3(new_n660), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n227), .A2(new_n228), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n230), .A2(new_n231), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n240), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n244), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n640), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n805), .A2(new_n811), .A3(KEYINPUT115), .A4(new_n660), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT116), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n814), .A2(new_n819), .A3(new_n823), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n814), .A2(new_n245), .A3(new_n820), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n667), .A2(new_n818), .A3(new_n669), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n696), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n799), .B1(new_n830), .B2(new_n614), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n580), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n534), .A2(new_n483), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n746), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT117), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n246), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n831), .A2(new_n534), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n580), .A2(new_n518), .A3(new_n521), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n482), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n246), .A2(new_n361), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  NOR3_X1   g642(.A1(new_n835), .A2(new_n371), .A3(new_n670), .ZN(new_n844));
  INV_X1    g643(.A(new_n841), .ZN(new_n845));
  AOI21_X1  g644(.A(G120gat), .B1(new_n845), .B2(new_n698), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(G1341gat));
  OAI21_X1  g646(.A(new_n381), .B1(new_n835), .B2(new_n614), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n614), .A2(new_n381), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n841), .B2(new_n849), .ZN(G1342gat));
  OAI21_X1  g649(.A(G134gat), .B1(new_n835), .B2(new_n696), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n845), .A2(new_n374), .A3(new_n376), .A4(new_n640), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n688), .A2(new_n833), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n580), .A2(KEYINPUT57), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n827), .B1(new_n246), .B2(new_n812), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n696), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(KEYINPUT119), .A3(new_n696), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n825), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n614), .ZN(new_n864));
  INV_X1    g663(.A(new_n799), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(new_n831), .B2(new_n581), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(KEYINPUT118), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n822), .A2(new_n824), .B1(new_n828), .B2(new_n696), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n865), .B1(new_n870), .B2(new_n699), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n580), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n856), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n254), .B1(new_n875), .B2(new_n245), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n726), .A2(new_n483), .A3(new_n581), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n837), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n246), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT58), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n856), .ZN(new_n881));
  INV_X1    g680(.A(new_n866), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n873), .B2(new_n872), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT118), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n245), .B(new_n881), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  INV_X1    g686(.A(new_n879), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n880), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(new_n878), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n256), .A3(new_n698), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n256), .C1(new_n875), .C2(new_n698), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n831), .B2(new_n581), .ZN(new_n895));
  INV_X1    g694(.A(new_n819), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(new_n812), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n699), .B1(new_n859), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n867), .B(new_n580), .C1(new_n898), .C2(new_n799), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n856), .A2(new_n670), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n256), .B1(new_n903), .B2(KEYINPUT121), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n900), .B2(new_n902), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n894), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n892), .B1(new_n893), .B2(new_n907), .ZN(G1345gat));
  AOI21_X1  g707(.A(KEYINPUT122), .B1(new_n891), .B2(new_n699), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n878), .A2(new_n910), .A3(new_n614), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n909), .A2(G155gat), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n614), .A2(new_n260), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n875), .B2(new_n913), .ZN(G1346gat));
  AOI21_X1  g713(.A(G162gat), .B1(new_n891), .B2(new_n640), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n696), .A2(new_n261), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n875), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n418), .A2(new_n482), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n832), .A2(new_n746), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(G169gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(new_n246), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n831), .A2(new_n418), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n483), .A3(new_n838), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(new_n246), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n924), .B2(new_n920), .ZN(G1348gat));
  OAI21_X1  g724(.A(G176gat), .B1(new_n919), .B2(new_n670), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n670), .A2(G176gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n923), .B2(new_n927), .ZN(G1349gat));
  OAI21_X1  g727(.A(G183gat), .B1(new_n919), .B2(new_n614), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n614), .A2(new_n437), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n919), .B2(new_n696), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n640), .A2(new_n428), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n934), .A2(new_n935), .B1(new_n923), .B2(new_n936), .ZN(G1351gat));
  NOR3_X1   g736(.A1(new_n726), .A2(new_n482), .A3(new_n581), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n245), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n895), .A2(new_n899), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n688), .A2(new_n918), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT123), .Z(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(G197gat), .A3(new_n245), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n941), .B1(new_n942), .B2(new_n945), .ZN(G1352gat));
  NOR3_X1   g745(.A1(new_n939), .A2(G204gat), .A3(new_n670), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n942), .A2(new_n698), .A3(new_n944), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n299), .B2(new_n949), .ZN(G1353gat));
  NAND2_X1  g749(.A1(new_n943), .A2(new_n699), .ZN(new_n951));
  OAI21_X1  g750(.A(G211gat), .B1(new_n900), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT63), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n954), .B(G211gat), .C1(new_n900), .C2(new_n951), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n614), .A2(G211gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n922), .A2(new_n938), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n938), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(new_n955), .A3(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n953), .A2(KEYINPUT125), .A3(new_n955), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1354gat));
  NAND2_X1  g765(.A1(new_n640), .A2(G218gat), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT126), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n942), .A2(new_n944), .A3(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G218gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n939), .B2(new_n696), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT127), .Z(G1355gat));
endmodule


