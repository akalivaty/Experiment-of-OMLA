

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n973), .ZN(n705) );
  NAND2_X1 U553 ( .A1(n798), .A2(n799), .ZN(n737) );
  XOR2_X1 U554 ( .A(KEYINPUT75), .B(n595), .Z(n973) );
  NAND2_X1 U555 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U556 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n719) );
  XNOR2_X1 U558 ( .A(n720), .B(n719), .ZN(n726) );
  NAND2_X1 U559 ( .A1(n726), .A2(n725), .ZN(n736) );
  INV_X1 U560 ( .A(KEYINPUT101), .ZN(n816) );
  XNOR2_X1 U561 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n591) );
  XNOR2_X1 U562 ( .A(n592), .B(n591), .ZN(n593) );
  NOR2_X1 U563 ( .A1(n641), .A2(n541), .ZN(n659) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n663) );
  INV_X1 U565 ( .A(KEYINPUT66), .ZN(n531) );
  XNOR2_X1 U566 ( .A(n532), .B(n531), .ZN(G160) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n521) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X2 U569 ( .A(n521), .B(n520), .ZN(n872) );
  NAND2_X1 U570 ( .A1(n872), .A2(G137), .ZN(n523) );
  INV_X1 U571 ( .A(G2105), .ZN(n526) );
  NOR2_X2 U572 ( .A1(G2104), .A2(n526), .ZN(n876) );
  NAND2_X1 U573 ( .A1(G125), .A2(n876), .ZN(n522) );
  AND2_X1 U574 ( .A1(n523), .A2(n522), .ZN(n530) );
  INV_X1 U575 ( .A(G2104), .ZN(n525) );
  NOR2_X4 U576 ( .A1(G2105), .A2(n525), .ZN(n871) );
  NAND2_X1 U577 ( .A1(G101), .A2(n871), .ZN(n524) );
  XNOR2_X1 U578 ( .A(KEYINPUT23), .B(n524), .ZN(n528) );
  NOR2_X2 U579 ( .A1(n526), .A2(n525), .ZN(n875) );
  AND2_X1 U580 ( .A1(n875), .A2(G113), .ZN(n527) );
  NOR2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U582 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n539) );
  XOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  NOR2_X1 U584 ( .A1(G651), .A2(n641), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT65), .B(n533), .Z(n655) );
  NAND2_X1 U586 ( .A1(n655), .A2(G51), .ZN(n537) );
  INV_X1 U587 ( .A(G651), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G543), .A2(n541), .ZN(n534) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n534), .Z(n535) );
  XNOR2_X1 U590 ( .A(KEYINPUT68), .B(n535), .ZN(n656) );
  NAND2_X1 U591 ( .A1(G63), .A2(n656), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n539), .B(n538), .ZN(n546) );
  NAND2_X1 U594 ( .A1(n663), .A2(G89), .ZN(n540) );
  XNOR2_X1 U595 ( .A(n540), .B(KEYINPUT4), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G76), .A2(n659), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U598 ( .A(KEYINPUT5), .B(n544), .Z(n545) );
  NOR2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U600 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n547) );
  XNOR2_X1 U601 ( .A(n548), .B(n547), .ZN(G168) );
  XOR2_X1 U602 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U603 ( .A1(n655), .A2(G47), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G60), .A2(n656), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G72), .A2(n659), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G85), .A2(n663), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U609 ( .A1(n554), .A2(n553), .ZN(G290) );
  XOR2_X1 U610 ( .A(G2430), .B(G2451), .Z(n556) );
  XNOR2_X1 U611 ( .A(KEYINPUT105), .B(G2443), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n556), .B(n555), .ZN(n563) );
  XOR2_X1 U613 ( .A(G2435), .B(G2446), .Z(n558) );
  XNOR2_X1 U614 ( .A(G2427), .B(G2454), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U616 ( .A(n559), .B(G2438), .Z(n561) );
  XNOR2_X1 U617 ( .A(G1341), .B(G1348), .ZN(n560) );
  XNOR2_X1 U618 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n563), .B(n562), .ZN(n564) );
  AND2_X1 U620 ( .A1(n564), .A2(G14), .ZN(G401) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  NAND2_X1 U625 ( .A1(n655), .A2(G52), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G64), .A2(n656), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G77), .A2(n659), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G90), .A2(n663), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U632 ( .A1(n571), .A2(n570), .ZN(G171) );
  INV_X1 U633 ( .A(G171), .ZN(G301) );
  NAND2_X1 U634 ( .A1(G114), .A2(n875), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G126), .A2(n876), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n579) );
  INV_X1 U637 ( .A(KEYINPUT89), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G102), .A2(n871), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G138), .A2(n872), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(G164) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n580) );
  XOR2_X1 U644 ( .A(n580), .B(KEYINPUT10), .Z(n922) );
  NAND2_X1 U645 ( .A1(n922), .A2(G567), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  NAND2_X1 U647 ( .A1(n655), .A2(G43), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT74), .B(n582), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n656), .A2(G56), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT14), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n594) );
  NAND2_X1 U652 ( .A1(n659), .A2(G68), .ZN(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT72), .B(n586), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n588) );
  NAND2_X1 U655 ( .A1(G81), .A2(n663), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n592) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U659 ( .A1(n973), .A2(G860), .ZN(G153) );
  NAND2_X1 U660 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U661 ( .A1(n656), .A2(G66), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT76), .ZN(n603) );
  NAND2_X1 U663 ( .A1(G54), .A2(n655), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G92), .A2(n663), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G79), .A2(n659), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT77), .B(n599), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT15), .B(n604), .ZN(n979) );
  INV_X1 U671 ( .A(n979), .ZN(n711) );
  INV_X1 U672 ( .A(G868), .ZN(n676) );
  NAND2_X1 U673 ( .A1(n711), .A2(n676), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G78), .A2(n659), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G91), .A2(n663), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G53), .A2(n655), .ZN(n609) );
  XOR2_X1 U679 ( .A(KEYINPUT69), .B(n609), .Z(n611) );
  NAND2_X1 U680 ( .A1(G65), .A2(n656), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n980) );
  XOR2_X1 U683 ( .A(n980), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U684 ( .A1(G299), .A2(G868), .ZN(n615) );
  NOR2_X1 U685 ( .A1(G286), .A2(n676), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT80), .B(n616), .ZN(G297) );
  INV_X1 U688 ( .A(G559), .ZN(n619) );
  NOR2_X1 U689 ( .A1(G860), .A2(n619), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n711), .A2(n617), .ZN(n618) );
  XOR2_X1 U691 ( .A(KEYINPUT16), .B(n618), .Z(G148) );
  NAND2_X1 U692 ( .A1(n619), .A2(n979), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n620), .A2(G868), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n705), .A2(n676), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G99), .A2(n871), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G111), .A2(n875), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n876), .A2(G123), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(KEYINPUT18), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G135), .A2(n872), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U703 ( .A(KEYINPUT81), .B(n628), .Z(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n929) );
  XNOR2_X1 U705 ( .A(G2096), .B(n929), .ZN(n631) );
  INV_X1 U706 ( .A(G2100), .ZN(n897) );
  NAND2_X1 U707 ( .A1(n631), .A2(n897), .ZN(G156) );
  NAND2_X1 U708 ( .A1(n655), .A2(G55), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G67), .A2(n656), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n659), .A2(G80), .ZN(n634) );
  XOR2_X1 U712 ( .A(KEYINPUT82), .B(n634), .Z(n635) );
  NOR2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n663), .A2(G93), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n675) );
  NAND2_X1 U716 ( .A1(n979), .A2(G559), .ZN(n673) );
  XOR2_X1 U717 ( .A(n973), .B(n673), .Z(n639) );
  NOR2_X1 U718 ( .A1(G860), .A2(n639), .ZN(n640) );
  XOR2_X1 U719 ( .A(n675), .B(n640), .Z(G145) );
  NAND2_X1 U720 ( .A1(G651), .A2(G74), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G49), .A2(n655), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G87), .A2(n641), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n656), .A2(n644), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(n647), .Z(G288) );
  NAND2_X1 U727 ( .A1(n655), .A2(G50), .ZN(n649) );
  NAND2_X1 U728 ( .A1(G62), .A2(n656), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U730 ( .A(KEYINPUT84), .B(n650), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G75), .A2(n659), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G88), .A2(n663), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U734 ( .A1(n654), .A2(n653), .ZN(G166) );
  NAND2_X1 U735 ( .A1(n655), .A2(G48), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G61), .A2(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n659), .A2(G73), .ZN(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n660), .Z(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n663), .A2(G86), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(G305) );
  XOR2_X1 U743 ( .A(G299), .B(n973), .Z(n672) );
  XOR2_X1 U744 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n666) );
  XNOR2_X1 U745 ( .A(G288), .B(n666), .ZN(n669) );
  XNOR2_X1 U746 ( .A(G166), .B(G305), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(n675), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n670), .B(G290), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n672), .B(n671), .ZN(n887) );
  XNOR2_X1 U751 ( .A(n673), .B(n887), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(G868), .ZN(n678) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U759 ( .A1(n682), .A2(G2072), .ZN(n683) );
  XNOR2_X1 U760 ( .A(KEYINPUT86), .B(n683), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U762 ( .A1(G120), .A2(G69), .ZN(n684) );
  NOR2_X1 U763 ( .A1(G237), .A2(n684), .ZN(n685) );
  XNOR2_X1 U764 ( .A(KEYINPUT88), .B(n685), .ZN(n686) );
  NAND2_X1 U765 ( .A1(n686), .A2(G108), .ZN(n842) );
  NAND2_X1 U766 ( .A1(n842), .A2(G567), .ZN(n692) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n687) );
  XNOR2_X1 U768 ( .A(KEYINPUT22), .B(n687), .ZN(n688) );
  NAND2_X1 U769 ( .A1(n688), .A2(G96), .ZN(n689) );
  NOR2_X1 U770 ( .A1(n689), .A2(G218), .ZN(n690) );
  XNOR2_X1 U771 ( .A(n690), .B(KEYINPUT87), .ZN(n843) );
  NAND2_X1 U772 ( .A1(n843), .A2(G2106), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n692), .A2(n691), .ZN(n921) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U775 ( .A1(n921), .A2(n693), .ZN(n841) );
  NAND2_X1 U776 ( .A1(n841), .A2(G36), .ZN(G176) );
  XOR2_X1 U777 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n694) );
  XNOR2_X1 U779 ( .A(n694), .B(KEYINPUT91), .ZN(n798) );
  NOR2_X1 U780 ( .A1(G1384), .A2(G164), .ZN(n695) );
  XNOR2_X1 U781 ( .A(n695), .B(KEYINPUT64), .ZN(n799) );
  AND2_X1 U782 ( .A1(n798), .A2(n799), .ZN(n722) );
  NAND2_X1 U783 ( .A1(n722), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U784 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  XNOR2_X1 U785 ( .A(G1956), .B(KEYINPUT97), .ZN(n1009) );
  NOR2_X1 U786 ( .A1(n1009), .A2(n722), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n714) );
  NOR2_X1 U788 ( .A1(n980), .A2(n714), .ZN(n700) );
  INV_X1 U789 ( .A(KEYINPUT28), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n700), .B(n699), .ZN(n718) );
  INV_X1 U791 ( .A(G1996), .ZN(n905) );
  NOR2_X1 U792 ( .A1(n737), .A2(n905), .ZN(n701) );
  XOR2_X1 U793 ( .A(n701), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U794 ( .A1(n737), .A2(G1341), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U797 ( .A1(G1348), .A2(n737), .ZN(n707) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n722), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n708) );
  OR2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n980), .A2(n714), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n722), .A2(G1961), .ZN(n721) );
  XOR2_X1 U807 ( .A(KEYINPUT96), .B(n721), .Z(n724) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n958) );
  NAND2_X1 U809 ( .A1(n722), .A2(n958), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n731) );
  NAND2_X1 U811 ( .A1(n731), .A2(G171), .ZN(n725) );
  NAND2_X1 U812 ( .A1(G8), .A2(n737), .ZN(n738) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n738), .ZN(n748) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n737), .ZN(n746) );
  NOR2_X1 U815 ( .A1(n748), .A2(n746), .ZN(n727) );
  XNOR2_X1 U816 ( .A(n727), .B(KEYINPUT98), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n728), .A2(G8), .ZN(n729) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n730), .A2(G168), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G171), .A2(n731), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n734), .Z(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n747) );
  NAND2_X1 U824 ( .A1(n747), .A2(G286), .ZN(n743) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n737), .ZN(n740) );
  BUF_X1 U826 ( .A(n738), .Z(n779) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n779), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U829 ( .A1(G303), .A2(n741), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(G8), .A2(n744), .ZN(n745) );
  XNOR2_X1 U832 ( .A(n745), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U833 ( .A1(G8), .A2(n746), .ZN(n751) );
  INV_X1 U834 ( .A(n747), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n753), .A2(n752), .ZN(n755) );
  INV_X1 U838 ( .A(KEYINPUT99), .ZN(n754) );
  XNOR2_X1 U839 ( .A(n755), .B(n754), .ZN(n773) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n758) );
  NOR2_X1 U841 ( .A1(G303), .A2(G1971), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n758), .A2(n756), .ZN(n996) );
  XOR2_X1 U843 ( .A(G1981), .B(KEYINPUT100), .Z(n757) );
  XNOR2_X1 U844 ( .A(G305), .B(n757), .ZN(n976) );
  INV_X1 U845 ( .A(n976), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n779), .A2(n759), .ZN(n760) );
  OR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n765) );
  INV_X1 U849 ( .A(n765), .ZN(n762) );
  AND2_X1 U850 ( .A1(n762), .A2(KEYINPUT33), .ZN(n768) );
  INV_X1 U851 ( .A(n768), .ZN(n763) );
  AND2_X1 U852 ( .A1(n996), .A2(n763), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n773), .A2(n764), .ZN(n770) );
  NOR2_X1 U854 ( .A1(n779), .A2(n765), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n984) );
  AND2_X1 U856 ( .A1(n766), .A2(n984), .ZN(n767) );
  OR2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n776) );
  NOR2_X1 U859 ( .A1(G303), .A2(G2090), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n774), .A2(n779), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U865 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n815) );
  NAND2_X1 U868 ( .A1(n875), .A2(G107), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G95), .A2(n871), .ZN(n782) );
  XOR2_X1 U870 ( .A(KEYINPUT93), .B(n782), .Z(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G119), .A2(n876), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G131), .A2(n872), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n851) );
  INV_X1 U876 ( .A(G1991), .ZN(n820) );
  NOR2_X1 U877 ( .A1(n851), .A2(n820), .ZN(n797) );
  NAND2_X1 U878 ( .A1(G117), .A2(n875), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G129), .A2(n876), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n871), .A2(G105), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n872), .A2(G141), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n867) );
  AND2_X1 U886 ( .A1(n867), .A2(G1996), .ZN(n796) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n927) );
  INV_X1 U888 ( .A(n798), .ZN(n800) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n833) );
  XOR2_X1 U890 ( .A(KEYINPUT94), .B(n833), .Z(n801) );
  NOR2_X1 U891 ( .A1(n927), .A2(n801), .ZN(n824) );
  INV_X1 U892 ( .A(n824), .ZN(n812) );
  NAND2_X1 U893 ( .A1(G104), .A2(n871), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G140), .A2(n872), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(KEYINPUT34), .B(n804), .ZN(n810) );
  NAND2_X1 U897 ( .A1(G116), .A2(n875), .ZN(n806) );
  NAND2_X1 U898 ( .A1(G128), .A2(n876), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U900 ( .A(KEYINPUT92), .B(n807), .Z(n808) );
  XNOR2_X1 U901 ( .A(KEYINPUT35), .B(n808), .ZN(n809) );
  NOR2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n811), .ZN(n884) );
  XNOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .ZN(n831) );
  NOR2_X1 U905 ( .A1(n884), .A2(n831), .ZN(n934) );
  NAND2_X1 U906 ( .A1(n833), .A2(n934), .ZN(n828) );
  NAND2_X1 U907 ( .A1(n812), .A2(n828), .ZN(n813) );
  XOR2_X1 U908 ( .A(KEYINPUT95), .B(n813), .Z(n814) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n817) );
  XNOR2_X1 U910 ( .A(n817), .B(n816), .ZN(n819) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U912 ( .A1(n985), .A2(n833), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n836) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n867), .ZN(n924) );
  AND2_X1 U915 ( .A1(n820), .A2(n851), .ZN(n930) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n821) );
  XNOR2_X1 U917 ( .A(KEYINPUT102), .B(n821), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n930), .A2(n822), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n924), .A2(n825), .ZN(n826) );
  XOR2_X1 U921 ( .A(KEYINPUT103), .B(n826), .Z(n827) );
  XNOR2_X1 U922 ( .A(KEYINPUT39), .B(n827), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n830), .B(KEYINPUT104), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n884), .A2(n831), .ZN(n939) );
  NAND2_X1 U926 ( .A1(n832), .A2(n939), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U929 ( .A(n837), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n922), .ZN(G217) );
  NAND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  XOR2_X1 U932 ( .A(KEYINPUT106), .B(n838), .Z(n839) );
  NAND2_X1 U933 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G108), .ZN(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  NAND2_X1 U943 ( .A1(G124), .A2(n876), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U945 ( .A1(n871), .A2(G100), .ZN(n845) );
  NAND2_X1 U946 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U947 ( .A1(G112), .A2(n875), .ZN(n848) );
  NAND2_X1 U948 ( .A1(G136), .A2(n872), .ZN(n847) );
  NAND2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U950 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U951 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n853) );
  XNOR2_X1 U952 ( .A(n851), .B(G162), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n866) );
  XNOR2_X1 U954 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n858) );
  NAND2_X1 U955 ( .A1(n871), .A2(G106), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT112), .ZN(n856) );
  NAND2_X1 U957 ( .A1(G142), .A2(n872), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n864) );
  NAND2_X1 U960 ( .A1(n876), .A2(G130), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n859), .B(KEYINPUT110), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G118), .A2(n875), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(KEYINPUT111), .B(n862), .Z(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n866), .B(n865), .Z(n869) );
  XOR2_X1 U967 ( .A(G164), .B(n867), .Z(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n929), .B(n870), .ZN(n883) );
  NAND2_X1 U970 ( .A1(G103), .A2(n871), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G139), .A2(n872), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n881) );
  NAND2_X1 U973 ( .A1(G115), .A2(n875), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G127), .A2(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n941) );
  XNOR2_X1 U978 ( .A(G160), .B(n941), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U981 ( .A1(G37), .A2(n886), .ZN(G395) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n887), .Z(n889) );
  XOR2_X1 U983 ( .A(G301), .B(G286), .Z(n888) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n890), .B(n979), .ZN(n891) );
  NOR2_X1 U986 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U987 ( .A(KEYINPUT42), .B(G2084), .Z(n893) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2078), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U990 ( .A(n894), .B(G2096), .Z(n896) );
  XNOR2_X1 U991 ( .A(G2090), .B(G2072), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n901) );
  XOR2_X1 U993 ( .A(KEYINPUT43), .B(G2678), .Z(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT107), .B(n897), .Z(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(n901), .B(n900), .Z(G227) );
  XOR2_X1 U997 ( .A(KEYINPUT108), .B(G1956), .Z(n903) );
  XNOR2_X1 U998 ( .A(G1986), .B(G1961), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n904), .B(KEYINPUT109), .Z(n907) );
  XOR2_X1 U1001 ( .A(n905), .B(G1991), .Z(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1003 ( .A(G1976), .B(G1981), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G1966), .B(G1971), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G2474), .B(KEYINPUT41), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(G229) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT116), .B(n914), .ZN(n920) );
  NOR2_X1 U1011 ( .A1(n921), .A2(G401), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n915), .B(KEYINPUT115), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n921), .ZN(G319) );
  INV_X1 U1019 ( .A(n922), .ZN(G223) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n950) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT119), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(n926), .B(KEYINPUT51), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n938) );
  XNOR2_X1 U1026 ( .A(G2084), .B(G160), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT117), .B(n931), .Z(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT118), .B(n936), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n947) );
  XOR2_X1 U1034 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n944), .Z(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(n945), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n948), .ZN(n949) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(n953), .B(KEYINPUT121), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G2072), .B(G33), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(n958), .B(G27), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G1996), .B(G32), .Z(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1057 ( .A(G2084), .B(KEYINPUT54), .Z(n966) );
  XNOR2_X1 U1058 ( .A(G34), .B(n966), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(n969), .Z(n971) );
  INV_X1 U1061 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n972), .ZN(n1030) );
  INV_X1 U1064 ( .A(G16), .ZN(n1026) );
  XOR2_X1 U1065 ( .A(n1026), .B(KEYINPUT56), .Z(n998) );
  NAND2_X1 U1066 ( .A1(G303), .A2(G1971), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n973), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n994) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(KEYINPUT57), .ZN(n992) );
  XNOR2_X1 U1072 ( .A(n979), .B(G1348), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1956), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n990) );
  XOR2_X1 U1075 ( .A(G1961), .B(G301), .Z(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT122), .ZN(n988) );
  INV_X1 U1077 ( .A(n984), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1028) );
  XOR2_X1 U1085 ( .A(G1986), .B(G24), .Z(n1001) );
  XNOR2_X1 U1086 ( .A(G22), .B(KEYINPUT127), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n999), .B(G1971), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT58), .B(n1004), .Z(n1023) );
  XOR2_X1 U1092 ( .A(G1961), .B(G5), .Z(n1017) );
  XOR2_X1 U1093 ( .A(G1341), .B(G19), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G6), .B(G1981), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT124), .B(n1008), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1009), .B(G20), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(KEYINPUT59), .B(G1348), .Z(n1012) );
  XNOR2_X1 U1101 ( .A(G4), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT60), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT125), .B(G1966), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G21), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(KEYINPUT126), .B(n1021), .Z(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

