//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT28), .Z(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AND2_X1   g006(.A1(KEYINPUT72), .A2(KEYINPUT26), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT72), .A2(KEYINPUT26), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n210), .B(KEYINPUT73), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n207), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(KEYINPUT71), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n205), .B(new_n206), .C1(new_n211), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n216), .A2(new_n217), .ZN(new_n223));
  NOR4_X1   g022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT68), .B(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n206), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n226), .A2(KEYINPUT69), .ZN(new_n227));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n206), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(KEYINPUT24), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(new_n226), .B2(KEYINPUT69), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n224), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n232), .B(KEYINPUT70), .Z(new_n233));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n223), .B1(new_n220), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n220), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n229), .A2(KEYINPUT64), .A3(KEYINPUT24), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n206), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n230), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT25), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n219), .B1(new_n233), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT74), .B1(new_n247), .B2(G120gat), .ZN(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G113gat), .ZN(new_n250));
  MUX2_X1   g049(.A(new_n248), .B(KEYINPUT74), .S(new_n250), .Z(new_n251));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(KEYINPUT75), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(KEYINPUT75), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n247), .A2(G120gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n254), .B1(new_n259), .B2(new_n250), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n253), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n246), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G227gat), .A2(G233gat), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT78), .B(KEYINPUT34), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n264), .B2(new_n265), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G15gat), .B(G43gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT77), .ZN(new_n272));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n263), .A2(G227gat), .A3(G233gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT76), .B(KEYINPUT33), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(KEYINPUT32), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n275), .B(KEYINPUT32), .C1(new_n274), .C2(new_n276), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n270), .A2(new_n279), .A3(new_n280), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT36), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT36), .ZN(new_n285));
  INV_X1    g084(.A(new_n283), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(new_n281), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT31), .B(G50gat), .Z(new_n289));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290));
  XOR2_X1   g089(.A(G211gat), .B(G218gat), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  INV_X1    g092(.A(G211gat), .ZN(new_n294));
  INV_X1    g093(.A(G218gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n292), .B(new_n293), .C1(KEYINPUT22), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(KEYINPUT22), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n291), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G155gat), .B(G162gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G141gat), .B(G148gat), .Z(new_n304));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305));
  AND2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT83), .B(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT2), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(new_n304), .A3(new_n301), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n300), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n297), .B1(new_n299), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT86), .B1(new_n298), .B2(new_n291), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n314), .B1(new_n322), .B2(new_n315), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n290), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n300), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n313), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(G228gat), .A3(G233gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n318), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(G22gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n330), .A2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n289), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n330), .A2(new_n332), .ZN(new_n337));
  INV_X1    g136(.A(new_n289), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n246), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n246), .A2(new_n317), .A3(new_n341), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n325), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n300), .A3(new_n343), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT37), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G8gat), .B(G36gat), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT79), .ZN(new_n351));
  XOR2_X1   g150(.A(G64gat), .B(G92gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(KEYINPUT37), .A3(new_n346), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT38), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n353), .B(KEYINPUT80), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT38), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n353), .B1(new_n345), .B2(new_n346), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n316), .A2(new_n365), .A3(new_n262), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n308), .A2(new_n258), .A3(new_n312), .A4(new_n261), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(KEYINPUT4), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(KEYINPUT84), .ZN(new_n370));
  OR3_X1    g169(.A1(new_n367), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT5), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(KEYINPUT85), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n316), .A2(new_n365), .A3(new_n262), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n367), .A2(KEYINPUT4), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n377), .B(new_n373), .C1(new_n369), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n313), .A2(new_n262), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n380), .A2(new_n367), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(KEYINPUT5), .C1(new_n373), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT85), .B1(new_n372), .B2(new_n375), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  AOI21_X1  g188(.A(KEYINPUT6), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n389), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n383), .B2(new_n384), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT6), .B(new_n391), .C1(new_n383), .C2(new_n384), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n355), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n358), .A2(new_n364), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n362), .A2(KEYINPUT30), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  AOI211_X1 g198(.A(new_n399), .B(new_n353), .C1(new_n345), .C2(new_n346), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n347), .A2(new_n359), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n373), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT39), .B(new_n403), .C1(new_n372), .C2(new_n373), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n389), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n372), .A2(KEYINPUT39), .A3(new_n373), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n407), .A2(KEYINPUT40), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(KEYINPUT40), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n392), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n340), .B1(new_n397), .B2(new_n412), .ZN(new_n413));
  OR3_X1    g212(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT81), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n394), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT81), .B1(new_n400), .B2(new_n401), .ZN(new_n416));
  INV_X1    g215(.A(new_n398), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n340), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n288), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  OR3_X1    g220(.A1(new_n286), .A2(new_n281), .A3(KEYINPUT88), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT35), .ZN(new_n423));
  AND4_X1   g222(.A1(new_n423), .A2(new_n402), .A3(new_n339), .A4(new_n336), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT88), .B1(new_n286), .B2(new_n281), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n422), .A2(new_n415), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n419), .A2(new_n282), .A3(new_n283), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT35), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G15gat), .B(G22gat), .ZN(new_n431));
  INV_X1    g230(.A(G1gat), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(KEYINPUT16), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  OAI21_X1  g234(.A(G8gat), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(G8gat), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n437), .B(new_n438), .C1(new_n432), .C2(new_n431), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n441));
  INV_X1    g240(.A(G57gat), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(G64gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(G64gat), .ZN(new_n444));
  INV_X1    g243(.A(G64gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(KEYINPUT97), .A3(G57gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n443), .A2(new_n446), .A3(KEYINPUT98), .A4(new_n444), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT9), .ZN(new_n452));
  OR3_X1    g251(.A1(new_n452), .A2(G71gat), .A3(G78gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(G71gat), .A2(G78gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457));
  AND3_X1   g256(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n445), .A2(G57gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n461), .A3(KEYINPUT95), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n452), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT95), .B1(new_n444), .B2(new_n461), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n457), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT95), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n445), .A2(G57gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n442), .A2(G64gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n462), .A3(new_n463), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n457), .B1(new_n472), .B2(new_n460), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n456), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT21), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n440), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT100), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G127gat), .B(G155gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n449), .A2(new_n450), .B1(new_n454), .B2(new_n453), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT96), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n466), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT99), .B1(new_n484), .B2(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g284(.A1(G231gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT99), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n474), .A2(new_n488), .A3(new_n475), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n487), .B1(new_n485), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n480), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n484), .A2(KEYINPUT99), .A3(KEYINPUT21), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n474), .B2(new_n475), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n485), .A2(new_n489), .A3(new_n487), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n479), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n492), .B2(new_n497), .ZN(new_n501));
  XOR2_X1   g300(.A(G183gat), .B(G211gat), .Z(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n490), .A2(new_n491), .A3(new_n480), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n479), .B1(new_n495), .B2(new_n496), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n498), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n478), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n500), .B2(new_n501), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n508), .A3(new_n502), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n477), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT14), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G36gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n524), .A3(KEYINPUT15), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n519), .ZN(new_n528));
  XOR2_X1   g327(.A(G43gat), .B(G50gat), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n520), .A2(new_n524), .A3(KEYINPUT15), .A4(new_n529), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(KEYINPUT17), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(G85gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n545), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT101), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n548), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT101), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n536), .A3(new_n551), .A4(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n533), .A2(new_n553), .B1(KEYINPUT41), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT102), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n562), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT103), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n561), .B(new_n563), .C1(new_n565), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n510), .A2(new_n513), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT104), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n510), .A2(KEYINPUT104), .A3(new_n513), .A4(new_n574), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n440), .A2(new_n531), .A3(KEYINPUT92), .A4(new_n532), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n436), .A2(new_n439), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n533), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n533), .A2(new_n582), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT13), .Z(new_n587));
  AND3_X1   g386(.A1(new_n585), .A2(KEYINPUT93), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT93), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(KEYINPUT90), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n440), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n535), .A2(new_n591), .A3(new_n536), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n533), .A2(new_n582), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT18), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n594), .A2(new_n595), .A3(new_n586), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n595), .A3(new_n586), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n597), .ZN(new_n601));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT11), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n216), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G197gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n590), .A2(new_n599), .A3(new_n601), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n587), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n585), .A2(KEYINPUT93), .A3(new_n587), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n610), .A2(new_n601), .A3(new_n611), .A4(new_n599), .ZN(new_n612));
  INV_X1    g411(.A(new_n606), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n474), .A2(new_n549), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n553), .B(new_n456), .C1(new_n467), .C2(new_n473), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n484), .A2(KEYINPUT10), .A3(new_n553), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(new_n619), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n624), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n430), .A2(new_n579), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n415), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n432), .ZN(G1324gat));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n402), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT42), .B1(new_n641), .B2(new_n438), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  MUX2_X1   g443(.A(KEYINPUT42), .B(new_n642), .S(new_n644), .Z(G1325gat));
  XNOR2_X1  g444(.A(new_n288), .B(KEYINPUT105), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G15gat), .B1(new_n638), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n422), .A2(new_n425), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(G15gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n638), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n638), .A2(new_n419), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  AOI21_X1  g453(.A(new_n574), .B1(new_n421), .B2(new_n429), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n510), .A2(new_n513), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n637), .ZN(new_n658));
  NOR4_X1   g457(.A1(new_n656), .A2(new_n415), .A3(new_n523), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n418), .A2(new_n419), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n364), .A2(new_n395), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n355), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT87), .B1(new_n355), .B2(KEYINPUT38), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n411), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n663), .B1(new_n668), .B2(new_n340), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n669), .A2(new_n288), .B1(new_n428), .B2(new_n426), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n662), .B1(new_n670), .B2(new_n574), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n655), .A2(KEYINPUT44), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n658), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n395), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n523), .B1(new_n675), .B2(new_n676), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n661), .B1(new_n677), .B2(new_n678), .ZN(G1328gat));
  NOR2_X1   g478(.A1(new_n656), .A2(new_n658), .ZN(new_n680));
  INV_X1    g479(.A(new_n402), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n515), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n674), .ZN(new_n684));
  OAI21_X1  g483(.A(G36gat), .B1(new_n684), .B2(new_n402), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1329gat));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n646), .A3(new_n674), .A4(new_n672), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(KEYINPUT108), .A3(G43gat), .ZN(new_n689));
  INV_X1    g488(.A(G43gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n649), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n680), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT108), .B1(new_n688), .B2(G43gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n288), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n673), .A2(new_n696), .A3(new_n674), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G43gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(KEYINPUT47), .A3(new_n692), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(G1330gat));
  NOR3_X1   g499(.A1(new_n656), .A2(new_n419), .A3(new_n658), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(G50gat), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n340), .A2(G50gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n684), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT48), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n702), .B(new_n706), .C1(new_n684), .C2(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1331gat));
  NAND3_X1  g507(.A1(new_n579), .A2(new_n616), .A3(new_n636), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n670), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n395), .B(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g512(.A(new_n402), .B(KEYINPUT110), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT111), .ZN(new_n717));
  OR2_X1    g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1333gat));
  NAND3_X1  g518(.A1(new_n710), .A2(G71gat), .A3(new_n646), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n710), .A2(KEYINPUT112), .A3(G71gat), .A4(new_n646), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n670), .A2(new_n649), .A3(new_n709), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n722), .B(new_n723), .C1(G71gat), .C2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n340), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G78gat), .ZN(G1335gat));
  INV_X1    g527(.A(new_n657), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n615), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n635), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n673), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n415), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n415), .A2(G85gat), .A3(new_n635), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n655), .A2(KEYINPUT113), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n730), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n655), .A2(KEYINPUT113), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n739), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n731), .B1(new_n655), .B2(KEYINPUT113), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT51), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n735), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(G1336gat));
  NOR3_X1   g544(.A1(new_n714), .A2(G92gat), .A3(new_n635), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n741), .A2(KEYINPUT51), .A3(new_n742), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n671), .A2(new_n681), .A3(new_n672), .A4(new_n732), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT52), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n746), .B1(new_n740), .B2(new_n743), .ZN(new_n754));
  INV_X1    g553(.A(new_n714), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n671), .A2(new_n672), .A3(new_n755), .A4(new_n732), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT52), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n758), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n733), .B2(new_n647), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n649), .A2(G99gat), .A3(new_n635), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n740), .B2(new_n743), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1338gat));
  NOR3_X1   g562(.A1(new_n419), .A2(G106gat), .A3(new_n635), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n748), .B2(new_n749), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n671), .A2(new_n340), .A3(new_n672), .A4(new_n732), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G106gat), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT53), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n740), .B2(new_n743), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(new_n768), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1339gat));
  NAND3_X1  g573(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n624), .A2(KEYINPUT54), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n626), .B1(new_n620), .B2(new_n621), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n633), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n607), .A2(new_n614), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(KEYINPUT55), .A3(new_n779), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n783), .A2(KEYINPUT114), .A3(new_n634), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT114), .B1(new_n783), .B2(new_n634), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n585), .A2(new_n587), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n605), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n607), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n635), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n573), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n780), .A2(new_n781), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n795), .A2(new_n573), .A3(new_n607), .A4(new_n790), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n783), .A2(new_n634), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT114), .A3(new_n634), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n794), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n800), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n574), .A2(new_n791), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n795), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n792), .B1(new_n804), .B2(new_n782), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n803), .B(new_n806), .C1(new_n807), .C2(new_n573), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n808), .A3(new_n657), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n577), .A2(new_n578), .A3(new_n616), .A4(new_n635), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n711), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n714), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n427), .ZN(new_n814));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n615), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n577), .A2(new_n578), .A3(new_n616), .A4(new_n635), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n786), .A2(new_n793), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n801), .B1(new_n817), .B2(new_n574), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n729), .B1(new_n818), .B2(new_n803), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n802), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n340), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n755), .A2(new_n415), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n691), .A3(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT116), .Z(new_n824));
  NOR2_X1   g623(.A1(new_n616), .A2(new_n247), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n815), .B1(new_n824), .B2(new_n825), .ZN(G1340gat));
  AOI21_X1  g625(.A(G120gat), .B1(new_n814), .B2(new_n636), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n635), .A2(new_n249), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n824), .B2(new_n828), .ZN(G1341gat));
  INV_X1    g628(.A(new_n824), .ZN(new_n830));
  OAI21_X1  g629(.A(G127gat), .B1(new_n830), .B2(new_n657), .ZN(new_n831));
  INV_X1    g630(.A(G127gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n832), .A3(new_n729), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1342gat));
  AND3_X1   g633(.A1(new_n812), .A2(new_n402), .A3(new_n573), .ZN(new_n835));
  INV_X1    g634(.A(G134gat), .ZN(new_n836));
  INV_X1    g635(.A(new_n427), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT117), .Z(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n830), .B2(new_n574), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n840), .B(new_n841), .C1(KEYINPUT56), .C2(new_n838), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n288), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n419), .B1(new_n809), .B2(new_n810), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(KEYINPUT57), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n782), .A2(new_n634), .A3(new_n783), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n573), .B1(new_n793), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n657), .B1(new_n848), .B2(new_n801), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n810), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n419), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n845), .A2(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT118), .B1(new_n844), .B2(KEYINPUT57), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n843), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(G141gat), .A3(new_n615), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n646), .A2(new_n419), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n714), .A3(new_n812), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n616), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(G141gat), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n846), .B(new_n851), .C1(new_n820), .C2(new_n419), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n850), .A2(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n854), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n843), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n636), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(G148gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(KEYINPUT59), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT119), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n810), .A2(KEYINPUT120), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n849), .B1(new_n810), .B2(KEYINPUT120), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n810), .A2(KEYINPUT120), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n849), .A4(new_n874), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n877), .A2(new_n879), .A3(new_n851), .A4(new_n340), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT57), .B1(new_n820), .B2(new_n419), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n636), .A3(new_n866), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n872), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n870), .A2(new_n871), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n858), .A2(G148gat), .A3(new_n635), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n862), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n885), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n882), .A2(G148gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT59), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n867), .A2(new_n869), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(KEYINPUT119), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT122), .B(new_n887), .C1(new_n891), .C2(new_n870), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n886), .A2(new_n892), .ZN(G1345gat));
  INV_X1    g692(.A(new_n855), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n657), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n729), .A2(new_n309), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n895), .A2(new_n309), .B1(new_n858), .B2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n894), .B2(new_n574), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n835), .A2(new_n310), .A3(new_n857), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  NAND2_X1  g699(.A1(new_n811), .A2(new_n415), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n837), .A3(new_n755), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n615), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n711), .A2(new_n402), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT124), .Z(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n691), .A3(new_n821), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n216), .A3(new_n616), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n905), .A2(new_n909), .ZN(G1348gat));
  OAI21_X1  g709(.A(G176gat), .B1(new_n908), .B2(new_n635), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n636), .A2(new_n217), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n903), .B2(new_n912), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n729), .A2(new_n202), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n903), .A2(KEYINPUT125), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n908), .B2(new_n657), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT125), .B1(new_n903), .B2(new_n914), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT60), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n915), .A2(new_n916), .A3(new_n920), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n908), .B2(new_n574), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n203), .A3(new_n573), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1351gat));
  XNOR2_X1  g726(.A(new_n906), .B(KEYINPUT124), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n646), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n880), .A2(new_n881), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n616), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n902), .A2(new_n755), .A3(new_n857), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n616), .A2(G197gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  INV_X1    g734(.A(G204gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n636), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n929), .A2(new_n636), .A3(new_n930), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n939), .A2(new_n940), .B1(new_n936), .B2(new_n941), .ZN(G1353gat));
  OAI21_X1  g741(.A(G211gat), .B1(new_n931), .B2(new_n657), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n729), .A2(new_n294), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n945), .A2(new_n946), .B1(new_n933), .B2(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(new_n295), .B1(new_n933), .B2(new_n574), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n929), .A2(new_n930), .A3(G218gat), .A4(new_n573), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(G1355gat));
endmodule


