//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n208), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n211), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  XOR2_X1   g0045(.A(KEYINPUT77), .B(KEYINPUT14), .Z(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  OAI211_X1 g0048(.A(G1), .B(G13), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n249), .A2(G274), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  AOI21_X1  g0051(.A(G1), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT74), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n249), .A2(G274), .ZN(new_n256));
  INV_X1    g0056(.A(new_n252), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT74), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n249), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n230), .A2(G1698), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G226), .B2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n264), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n249), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n263), .A2(G238), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n260), .A2(new_n261), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n260), .B2(new_n273), .ZN(new_n276));
  OAI211_X1 g0076(.A(G169), .B(new_n246), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n260), .A2(new_n273), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n274), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n277), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n280), .B2(new_n274), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT76), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(G169), .B1(new_n275), .B2(new_n276), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT76), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT14), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n282), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n206), .A3(G1), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT12), .B1(new_n293), .B2(G68), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n224), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G68), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n205), .B2(G20), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n294), .A2(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G50), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n247), .A2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n308), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n297), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n301), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n290), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n275), .A2(new_n276), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(G190), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT75), .B1(new_n281), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n314), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT17), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n205), .A2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n298), .B1(new_n292), .B2(new_n330), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT79), .ZN(new_n336));
  INV_X1    g0136(.A(new_n297), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT7), .B1(new_n270), .B2(new_n206), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n339), .B(G20), .C1(new_n268), .C2(new_n269), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G58), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n299), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G58), .A2(G68), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n302), .A2(new_n303), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(G20), .B1(new_n346), .B2(G159), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n337), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n247), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT3), .B(G33), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(KEYINPUT78), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n339), .B1(new_n353), .B2(new_n206), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT78), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT78), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(new_n267), .A3(G33), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n355), .A2(new_n339), .A3(new_n206), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G68), .ZN(new_n359));
  OAI211_X1 g0159(.A(KEYINPUT16), .B(new_n347), .C1(new_n354), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n336), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n339), .B1(new_n352), .B2(G20), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n299), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n343), .B2(new_n344), .ZN(new_n365));
  INV_X1    g0165(.A(G159), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n304), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n349), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  AND4_X1   g0168(.A1(new_n336), .A2(new_n360), .A3(new_n297), .A4(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n335), .B1(new_n361), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G226), .A2(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT80), .B1(new_n353), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(new_n357), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT80), .ZN(new_n374));
  INV_X1    g0174(.A(new_n371), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G87), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n247), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G1698), .B1(new_n355), .B2(new_n357), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(G223), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n249), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n253), .B1(new_n230), .B2(new_n262), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n323), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n353), .A2(KEYINPUT80), .A3(new_n371), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n374), .B1(new_n373), .B2(new_n375), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n272), .ZN(new_n388));
  INV_X1    g0188(.A(new_n383), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n320), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n329), .B1(new_n370), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n335), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n360), .A2(new_n368), .A3(new_n297), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT79), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n350), .A2(new_n336), .A3(new_n360), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n283), .B1(new_n388), .B2(new_n389), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n278), .B(new_n383), .C1(new_n387), .C2(new_n272), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n382), .B2(new_n383), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n388), .A2(new_n389), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n278), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n370), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n384), .A2(new_n390), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n392), .A2(new_n401), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n298), .A2(G77), .A3(new_n332), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT71), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n202), .B2(new_n292), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n308), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT69), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n346), .A2(new_n331), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G20), .A2(G77), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT70), .A3(new_n297), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT70), .B1(new_n420), .B2(new_n297), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n413), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n258), .B1(G244), .B2(new_n263), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n352), .A2(G1698), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT66), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G238), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n270), .A2(new_n230), .A3(G1698), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT68), .B(G107), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n270), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n278), .B(new_n425), .C1(new_n432), .C2(new_n249), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n249), .B1(new_n428), .B2(new_n431), .ZN(new_n434));
  INV_X1    g0234(.A(new_n425), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n283), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n424), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n258), .B1(G226), .B2(new_n263), .ZN(new_n438));
  INV_X1    g0238(.A(G1698), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n352), .A2(G222), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n202), .B2(new_n352), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n427), .B2(G223), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n438), .B1(new_n442), .B2(new_n249), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n283), .ZN(new_n444));
  INV_X1    g0244(.A(G150), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n304), .A2(new_n445), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n330), .A2(new_n308), .B1(new_n206), .B2(new_n201), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n297), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n305), .B1(new_n205), .B2(G20), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n298), .A2(new_n449), .B1(new_n305), .B2(new_n292), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n444), .B(new_n451), .C1(G179), .C2(new_n443), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n420), .A2(new_n297), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT70), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n421), .ZN(new_n456));
  OAI211_X1 g0256(.A(G190), .B(new_n425), .C1(new_n432), .C2(new_n249), .ZN(new_n457));
  OAI21_X1  g0257(.A(G200), .B1(new_n434), .B2(new_n435), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n413), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n437), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT10), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n461), .A2(KEYINPUT10), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT72), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n443), .A2(new_n464), .A3(G200), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n451), .B(KEYINPUT9), .ZN(new_n466));
  OAI211_X1 g0266(.A(G190), .B(new_n438), .C1(new_n442), .C2(new_n249), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n464), .B1(new_n443), .B2(G200), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n462), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n468), .ZN(new_n471));
  INV_X1    g0271(.A(new_n469), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n471), .A2(new_n461), .A3(KEYINPUT10), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n460), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n328), .A2(new_n410), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n292), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n298), .B1(G1), .B2(new_n247), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n477), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT6), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n482), .A2(new_n477), .A3(G107), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(G20), .B1(G77), .B2(new_n346), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n430), .B1(new_n338), .B2(new_n340), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n480), .B1(new_n489), .B2(new_n297), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n213), .B1(new_n355), .B2(new_n357), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT4), .B1(new_n491), .B2(new_n439), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n493), .A2(new_n213), .A3(G1698), .ZN(new_n494));
  INV_X1    g0294(.A(G250), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n439), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n352), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n272), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n205), .A2(G45), .ZN(new_n501));
  OR2_X1    g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n504), .A2(G274), .A3(new_n249), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n272), .A2(new_n504), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(G257), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n500), .A2(G190), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n490), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n323), .B1(new_n500), .B2(new_n507), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT81), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n510), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT81), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n490), .A4(new_n508), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n414), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n293), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(new_n297), .B(new_n292), .C1(new_n205), .C2(G33), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n516), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT19), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n307), .A2(new_n521), .A3(G97), .ZN(new_n522));
  AND2_X1   g0322(.A1(KEYINPUT68), .A2(G107), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT68), .A2(G107), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G87), .A2(G97), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(new_n206), .B2(new_n264), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n522), .B1(new_n527), .B2(new_n521), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n373), .A2(new_n206), .A3(G68), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n518), .B(new_n520), .C1(new_n530), .C2(new_n337), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n380), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n491), .A2(G1698), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n249), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n501), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n249), .A2(G274), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n249), .A2(G250), .A3(new_n501), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT82), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT82), .B1(new_n537), .B2(new_n536), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n283), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n373), .A2(G238), .A3(new_n439), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n533), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n272), .ZN(new_n546));
  INV_X1    g0346(.A(new_n540), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n538), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n278), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n531), .A2(new_n542), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(G200), .B1(new_n534), .B2(new_n541), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(G190), .A3(new_n548), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n337), .B1(new_n528), .B2(new_n529), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n479), .A2(new_n378), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n553), .A2(new_n517), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n500), .A2(new_n278), .A3(new_n507), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n484), .B1(new_n482), .B2(new_n481), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n559), .A2(new_n206), .B1(new_n304), .B2(new_n202), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n525), .B1(new_n362), .B2(new_n363), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n297), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n519), .A2(G97), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n478), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n506), .A2(G257), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n250), .A2(new_n504), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n499), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n353), .A2(new_n213), .A3(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(KEYINPUT4), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n570), .B2(new_n272), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n558), .B(new_n564), .C1(new_n571), .C2(G169), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n515), .A2(new_n557), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n292), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n479), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n498), .B(new_n206), .C1(G33), .C2(new_n477), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT83), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n296), .A2(new_n224), .B1(G20), .B2(new_n575), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n578), .A2(KEYINPUT83), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  AOI21_X1  g0385(.A(G20), .B1(G33), .B2(G283), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n247), .A2(G97), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT20), .B(new_n580), .C1(new_n584), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n577), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n506), .A2(G270), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G257), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n215), .B2(G1698), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n373), .A2(new_n593), .B1(G303), .B2(new_n270), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n591), .B(new_n566), .C1(new_n594), .C2(new_n249), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G169), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n574), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n519), .A2(G116), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT20), .B1(new_n579), .B2(new_n580), .ZN(new_n599));
  INV_X1    g0399(.A(new_n589), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n576), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n595), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(G179), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n601), .A2(KEYINPUT21), .A3(G169), .A4(new_n595), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(G190), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(G200), .B2(new_n595), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT23), .B1(new_n430), .B2(new_n206), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n430), .C2(new_n206), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT23), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n206), .A2(G107), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n307), .B2(G116), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n206), .A2(G87), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n270), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI211_X1 g0423(.A(G20), .B(new_n378), .C1(new_n355), .C2(new_n357), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT22), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n610), .B1(new_n619), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n373), .A2(new_n206), .A3(G87), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n628), .B2(KEYINPUT22), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n629), .A2(new_n618), .A3(KEYINPUT24), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n297), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n291), .A2(G1), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT86), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(new_n616), .C1(new_n633), .C2(KEYINPUT25), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT25), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n519), .A2(G107), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n506), .A2(G264), .B1(new_n250), .B2(new_n504), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n495), .A2(new_n439), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(G257), .B2(new_n439), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n357), .B2(new_n355), .ZN(new_n643));
  INV_X1    g0443(.A(G294), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n247), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n272), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT87), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(new_n646), .A3(KEYINPUT87), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G169), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n640), .A2(new_n646), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G179), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n639), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(G190), .B1(new_n649), .B2(new_n650), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n652), .A2(G200), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n631), .B(new_n638), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NOR4_X1   g0459(.A1(new_n476), .A2(new_n573), .A3(new_n609), .A4(new_n659), .ZN(G372));
  AOI21_X1  g0460(.A(new_n324), .B1(new_n319), .B2(new_n321), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n437), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n315), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n392), .A2(new_n408), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n401), .A2(new_n406), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n473), .A2(KEYINPUT88), .A3(new_n470), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT88), .B1(new_n473), .B2(new_n470), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n452), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n550), .A2(new_n556), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n572), .ZN(new_n673));
  INV_X1    g0473(.A(new_n572), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(KEYINPUT26), .A3(new_n550), .A4(new_n556), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n550), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n631), .A2(new_n638), .B1(new_n651), .B2(new_n653), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n658), .B1(new_n678), .B2(new_n605), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n573), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n670), .B1(new_n476), .B2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n632), .A2(new_n206), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n659), .B1(new_n639), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT90), .Z(new_n690));
  NAND2_X1  g0490(.A1(new_n678), .A2(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n688), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n590), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n605), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n609), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT89), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n605), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n688), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n690), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n678), .A2(new_n694), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n209), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n525), .A2(new_n575), .A3(new_n526), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n205), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n223), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  OAI21_X1  g0514(.A(new_n591), .B1(new_n594), .B2(new_n249), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n647), .A2(new_n715), .A3(new_n278), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n534), .A2(new_n541), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n571), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n602), .A2(new_n652), .A3(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n500), .A2(new_n507), .ZN(new_n722));
  INV_X1    g0522(.A(new_n717), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT30), .A4(new_n571), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n688), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n727), .B(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT91), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n608), .A2(new_n655), .A3(new_n658), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n674), .B1(new_n511), .B2(new_n514), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n557), .A4(new_n694), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n729), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n702), .A2(new_n655), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(new_n735), .A3(new_n557), .A4(new_n658), .ZN(new_n740));
  INV_X1    g0540(.A(new_n550), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n673), .B2(new_n675), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n688), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n714), .B1(new_n746), .B2(G1), .ZN(G364));
  XOR2_X1   g0547(.A(new_n699), .B(KEYINPUT92), .Z(new_n748));
  NOR2_X1   g0548(.A1(new_n291), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n205), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n710), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n748), .B(new_n753), .C1(G330), .C2(new_n698), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n709), .A2(new_n270), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G355), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G116), .B2(new_n209), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n709), .A2(new_n373), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n251), .B2(new_n223), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n244), .A2(G45), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(G20), .B1(KEYINPUT93), .B2(G169), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(KEYINPUT93), .A2(G169), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n224), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n752), .B1(new_n762), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT95), .B1(new_n320), .B2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n320), .A2(KEYINPUT95), .A3(G20), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n323), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT97), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G283), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n206), .A2(new_n320), .A3(new_n323), .A4(G179), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n352), .B1(new_n780), .B2(G303), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n206), .A2(new_n278), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n320), .A3(new_n323), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI221_X1 g0588(.A(new_n781), .B1(new_n782), .B2(new_n784), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n320), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT94), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n789), .B1(G322), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n785), .A2(new_n320), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n790), .A2(new_n278), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(G326), .B1(new_n801), .B2(G294), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT98), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n776), .A2(G200), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n802), .A2(KEYINPUT98), .B1(new_n804), .B2(G329), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n779), .A2(new_n798), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n778), .A2(G107), .ZN(new_n807));
  INV_X1    g0607(.A(new_n801), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n477), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n787), .A2(new_n299), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(G50), .C2(new_n799), .ZN(new_n811));
  INV_X1    g0611(.A(new_n780), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n352), .B1(new_n202), .B2(new_n784), .C1(new_n812), .C2(new_n378), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n797), .B2(G58), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n807), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n804), .A2(G159), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n806), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n772), .B1(new_n819), .B2(new_n766), .ZN(new_n820));
  INV_X1    g0620(.A(new_n769), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n697), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n754), .A2(new_n822), .ZN(G396));
  AND4_X1   g0623(.A1(new_n424), .A2(new_n433), .A3(new_n436), .A4(new_n694), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n424), .A2(new_n688), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n459), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n824), .B1(new_n826), .B2(new_n437), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n827), .B(new_n694), .C1(new_n677), .C2(new_n680), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT101), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n743), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n743), .B2(new_n827), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n752), .B1(new_n833), .B2(new_n738), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n738), .B2(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n778), .A2(G87), .ZN(new_n836));
  INV_X1    g0636(.A(new_n799), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n809), .B(new_n839), .C1(G283), .C2(new_n786), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n270), .B1(new_n575), .B2(new_n784), .C1(new_n812), .C2(new_n214), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n797), .B2(G294), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n804), .A2(G311), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n836), .A2(new_n840), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n778), .A2(G68), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n373), .B1(new_n812), .B2(new_n305), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G58), .B2(new_n801), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  INV_X1    g0648(.A(new_n804), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n845), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n784), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G137), .A2(new_n799), .B1(new_n851), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n445), .B2(new_n787), .C1(new_n796), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n766), .ZN(new_n858));
  INV_X1    g0658(.A(new_n766), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n768), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n753), .B1(new_n862), .B2(new_n202), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n858), .B(new_n863), .C1(new_n827), .C2(new_n768), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n835), .A2(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n749), .A2(new_n205), .ZN(new_n866));
  INV_X1    g0666(.A(G330), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n736), .A2(new_n728), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n826), .A2(new_n437), .ZN(new_n869));
  INV_X1    g0669(.A(new_n824), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n314), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n688), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n326), .B(new_n873), .C1(new_n290), .C2(new_n314), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n284), .A2(new_n246), .B1(new_n317), .B2(G179), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n284), .A2(KEYINPUT76), .A3(new_n285), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n288), .B1(new_n287), .B2(KEYINPUT14), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n872), .B(new_n688), .C1(new_n878), .C2(new_n661), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n871), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n868), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n360), .A2(new_n297), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n347), .B1(new_n354), .B2(new_n359), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n349), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n393), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n686), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n409), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n409), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n397), .A2(new_n407), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n886), .B1(new_n400), .B2(new_n686), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n370), .A2(new_n405), .ZN(new_n897));
  INV_X1    g0697(.A(new_n686), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n370), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n897), .A2(new_n899), .A3(new_n893), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n892), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n409), .A2(new_n890), .A3(new_n887), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n890), .B1(new_n409), .B2(new_n887), .ZN(new_n905));
  OAI211_X1 g0705(.A(KEYINPUT38), .B(new_n902), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n882), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n881), .B1(new_n914), .B2(new_n906), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT105), .B1(new_n915), .B2(KEYINPUT40), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n897), .A2(new_n899), .A3(new_n893), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n901), .ZN(new_n920));
  INV_X1    g0720(.A(new_n899), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n409), .A2(KEYINPUT103), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT103), .B1(new_n409), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n906), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n868), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT106), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n476), .B1(new_n728), .B2(new_n736), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n867), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n476), .A2(new_n744), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n670), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT104), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT39), .B1(new_n925), .B2(new_n906), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n903), .A2(new_n907), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n938), .B2(KEYINPUT39), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n316), .A2(new_n688), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n938), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n829), .A2(new_n831), .A3(new_n870), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n874), .A2(new_n879), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n942), .A2(new_n946), .B1(new_n666), .B2(new_n686), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n936), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n866), .B1(new_n933), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n933), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(G116), .A3(new_n225), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n223), .B(G77), .C1(new_n342), .C2(new_n299), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(G50), .B2(new_n299), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(G1), .A3(new_n291), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(G367));
  OAI221_X1 g0759(.A(new_n770), .B1(new_n209), .B2(new_n414), .C1(new_n759), .C2(new_n236), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT109), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n753), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n808), .A2(new_n299), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n837), .A2(new_n853), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(G159), .C2(new_n786), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n352), .B1(new_n784), .B2(new_n305), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G58), .B2(new_n780), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(new_n445), .C2(new_n796), .ZN(new_n969));
  INV_X1    g0769(.A(new_n777), .ZN(new_n970));
  INV_X1    g0770(.A(G137), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n202), .A2(new_n970), .B1(new_n849), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT46), .B1(new_n780), .B2(G116), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n837), .B2(new_n782), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(G317), .C2(new_n804), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n477), .B2(new_n970), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n786), .A2(G294), .B1(new_n801), .B2(new_n430), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n373), .B1(G283), .B2(new_n851), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n796), .C2(new_n838), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n969), .A2(new_n972), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n963), .B1(new_n982), .B2(new_n766), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n555), .A2(new_n694), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n741), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n672), .B2(new_n984), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(new_n821), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n750), .B(KEYINPUT108), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n705), .A2(new_n706), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n735), .B1(new_n490), .B2(new_n694), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n674), .A2(new_n688), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n707), .A2(new_n994), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT45), .B1(new_n707), .B2(new_n994), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n700), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n999), .B(new_n1000), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n701), .A3(new_n998), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n705), .B1(new_n692), .B2(new_n703), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n748), .A2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n699), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n746), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1004), .A2(new_n1006), .A3(new_n1011), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1012), .A2(new_n746), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n710), .B(KEYINPUT41), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n990), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n705), .A2(new_n995), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT42), .Z(new_n1017));
  OAI21_X1  g0817(.A(new_n572), .B1(new_n992), .B2(new_n655), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(new_n694), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT107), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n986), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n701), .A2(new_n995), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n989), .B1(new_n1015), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n745), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n710), .A3(new_n1010), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n990), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1008), .A2(new_n1009), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n786), .B1(new_n851), .B2(G303), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n799), .A2(G322), .ZN(new_n1038));
  INV_X1    g0838(.A(G317), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1038), .C1(new_n796), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n801), .A2(G283), .B1(new_n780), .B2(G294), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT49), .Z(new_n1046));
  AOI21_X1  g0846(.A(new_n373), .B1(new_n804), .B2(G326), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n575), .B2(new_n970), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n808), .A2(new_n414), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n797), .B2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n799), .A2(G159), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT113), .Z(new_n1054));
  NOR2_X1   g0854(.A1(new_n787), .A2(new_n330), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n373), .B1(new_n299), .B2(new_n784), .C1(new_n812), .C2(new_n202), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n445), .B2(new_n849), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1052), .B(new_n1058), .C1(G97), .C2(new_n778), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1049), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n711), .A2(KEYINPUT110), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n711), .A2(KEYINPUT110), .ZN(new_n1062));
  AOI21_X1  g0862(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT111), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT111), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n330), .A2(G50), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT50), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n758), .C1(new_n251), .C2(new_n233), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n755), .A2(new_n711), .B1(new_n214), .B2(new_n709), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n752), .B1(new_n1072), .B2(new_n771), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1060), .A2(new_n766), .B1(KEYINPUT112), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(KEYINPUT112), .B2(new_n1073), .C1(new_n692), .C2(new_n821), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1036), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1034), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1034), .A2(KEYINPUT115), .A3(new_n1076), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(G393));
  NAND2_X1  g0881(.A1(new_n1012), .A2(new_n710), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1005), .A2(new_n701), .A3(new_n998), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n701), .B1(new_n1005), .B2(new_n998), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1010), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(KEYINPUT117), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT117), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n1010), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1004), .A2(new_n1006), .A3(new_n1035), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n241), .A2(new_n758), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n770), .B1(new_n477), .B2(new_n209), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n752), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n797), .A2(G311), .B1(G317), .B2(new_n799), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n787), .A2(new_n838), .B1(new_n808), .B2(new_n575), .ZN(new_n1100));
  INV_X1    g0900(.A(G283), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n270), .B1(new_n644), .B2(new_n784), .C1(new_n812), .C2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G322), .C2(new_n804), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1098), .A2(new_n807), .A3(new_n1099), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n796), .A2(new_n366), .B1(new_n445), .B2(new_n837), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT51), .Z(new_n1106));
  NAND2_X1  g0906(.A1(new_n804), .A2(G143), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n812), .A2(new_n299), .B1(new_n330), .B2(new_n784), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n353), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n808), .A2(new_n202), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G50), .B2(new_n786), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n836), .A2(new_n1107), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1104), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1095), .B1(new_n1113), .B2(new_n766), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n994), .B2(new_n821), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1092), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1091), .A2(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(new_n710), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n867), .B1(new_n736), .B2(new_n728), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n880), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT39), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n926), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n940), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1124), .A2(new_n1125), .B1(new_n945), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n828), .A2(new_n870), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n940), .B1(new_n1128), .B2(new_n944), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n926), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1122), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n737), .A2(G330), .A3(new_n827), .A4(new_n944), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1130), .B(new_n1133), .C1(new_n939), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1120), .A2(new_n827), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n944), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1128), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1133), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n737), .A2(G330), .A3(new_n827), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1122), .B1(new_n1142), .B2(new_n1139), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n943), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1120), .A2(new_n328), .A3(new_n410), .A4(new_n475), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n670), .A2(new_n934), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT118), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1119), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n939), .A2(new_n768), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n804), .A2(G125), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n352), .C1(new_n970), .C2(new_n305), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT119), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n799), .A2(G128), .B1(new_n801), .B2(G159), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n780), .A2(G150), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT53), .Z(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n787), .A2(new_n971), .B1(new_n784), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n797), .B2(G132), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n787), .A2(new_n525), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1110), .B(new_n1164), .C1(G283), .C2(new_n799), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n270), .B1(new_n477), .B2(new_n784), .C1(new_n812), .C2(new_n378), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n797), .B2(G116), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n804), .A2(G294), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n845), .A2(new_n1165), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n859), .B1(new_n1163), .B2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n753), .B(new_n1170), .C1(new_n330), .C2(new_n862), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT120), .Z(new_n1172));
  AOI22_X1  g0972(.A1(new_n1137), .A2(new_n1035), .B1(new_n1153), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1152), .A2(new_n1173), .ZN(G378));
  INV_X1    g0974(.A(KEYINPUT124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n452), .B1(new_n667), .B2(new_n668), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n451), .A2(new_n898), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n452), .B(new_n1177), .C1(new_n667), .C2(new_n668), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n928), .A2(G330), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n917), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1186), .B(new_n1188), .C1(new_n911), .C2(new_n916), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT123), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1190), .A2(new_n1191), .B1(new_n948), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n915), .A2(KEYINPUT105), .A3(KEYINPUT40), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1186), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1192), .B1(new_n941), .B2(new_n947), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n917), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n990), .B1(new_n1193), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n752), .B1(G50), .B2(new_n860), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n247), .A2(new_n248), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G50), .B(new_n1204), .C1(new_n248), .C2(new_n353), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G41), .B(new_n373), .C1(new_n797), .C2(G107), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n787), .A2(new_n477), .B1(new_n837), .B2(new_n575), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n812), .A2(new_n202), .B1(new_n414), .B2(new_n784), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1207), .A2(new_n964), .A3(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G58), .A2(new_n777), .B1(new_n804), .B2(G283), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1205), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n812), .A2(new_n1160), .B1(new_n784), .B2(new_n971), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G132), .B2(new_n786), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n799), .A2(G125), .B1(new_n801), .B2(G150), .ZN(new_n1216));
  INV_X1    g1016(.A(G128), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1215), .B(new_n1216), .C1(new_n1217), .C2(new_n796), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n777), .A2(G159), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n804), .A2(G124), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1204), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1202), .B1(new_n1224), .B2(new_n766), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1186), .B2(new_n768), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT122), .Z(new_n1227));
  OAI21_X1  g1027(.A(new_n1175), .B1(new_n1201), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1198), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1035), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1227), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT124), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n941), .A2(new_n947), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1197), .A2(new_n948), .A3(new_n1199), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1132), .A2(new_n1135), .A3(new_n1145), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1148), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT57), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1234), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1239), .B2(new_n1148), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1244), .A2(new_n1236), .A3(KEYINPUT125), .A4(new_n1237), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1193), .A2(new_n1200), .B1(new_n1148), .B2(new_n1239), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n710), .B1(new_n1247), .B2(KEYINPUT57), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1228), .B(new_n1233), .C1(new_n1246), .C2(new_n1248), .ZN(G375));
  OR2_X1    g1049(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1014), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1149), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1139), .A2(new_n767), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n752), .B1(new_n861), .B2(G68), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1050), .B1(G116), .B2(new_n786), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n644), .B2(new_n837), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n796), .A2(new_n1101), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n270), .B1(new_n525), .B2(new_n784), .C1(new_n812), .C2(new_n477), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n838), .B2(new_n849), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n778), .A2(G77), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n812), .A2(new_n366), .B1(new_n784), .B2(new_n445), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n353), .B(new_n1262), .C1(new_n797), .C2(G137), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n799), .A2(G132), .B1(new_n801), .B2(G50), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n787), .C2(new_n1160), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n342), .A2(new_n970), .B1(new_n849), .B2(new_n1217), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1260), .A2(new_n1261), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1254), .B1(new_n1267), .B2(new_n766), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1145), .A2(new_n1035), .B1(new_n1253), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1252), .A2(new_n1269), .ZN(G381));
  NOR2_X1   g1070(.A1(G390), .A2(G384), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  INV_X1    g1072(.A(G396), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1079), .A2(new_n1273), .A3(new_n1080), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G381), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1271), .A2(new_n1030), .A3(new_n1272), .A4(new_n1275), .ZN(G407));
  INV_X1    g1076(.A(G213), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(G343), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1272), .A2(new_n1278), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT126), .Z(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1081(.A(new_n1274), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1273), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1091), .B(new_n1117), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1086), .A2(KEYINPUT117), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1089), .A2(new_n1088), .A3(new_n1010), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1082), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1285), .B(new_n1274), .C1(new_n1288), .C2(new_n1116), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1284), .A2(new_n1289), .A3(new_n1030), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1030), .B1(new_n1284), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1236), .A2(new_n1237), .A3(new_n1035), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1152), .A2(new_n1173), .A3(new_n1232), .A4(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1240), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(new_n1014), .ZN(new_n1296));
  OAI22_X1  g1096(.A1(new_n1294), .A2(new_n1296), .B1(new_n1277), .B2(G343), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(G378), .B2(G375), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1299), .A2(new_n1250), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n710), .B1(new_n1299), .B2(new_n1250), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1269), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n835), .A3(new_n864), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G384), .B(new_n1269), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1233), .A2(new_n1228), .ZN(new_n1309));
  OAI21_X1  g1109(.A(G378), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1297), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1306), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1278), .A2(G2897), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1305), .B(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1292), .A2(new_n1307), .A3(new_n1314), .A4(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT62), .B1(new_n1298), .B2(new_n1306), .ZN(new_n1320));
  INV_X1    g1120(.A(G378), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1233), .A2(new_n1228), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1295), .A2(new_n1243), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1323), .A2(new_n710), .A3(new_n1242), .A4(new_n1245), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1321), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(new_n1325), .A2(new_n1326), .A3(new_n1305), .A4(new_n1297), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1318), .B(KEYINPUT127), .C1(new_n1320), .C2(new_n1327), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1312), .A2(new_n1326), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1298), .A2(KEYINPUT62), .A3(new_n1306), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT127), .B1(new_n1333), .B2(new_n1318), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1319), .B1(new_n1330), .B2(new_n1334), .ZN(G405));
  NOR2_X1   g1135(.A1(new_n1272), .A2(new_n1325), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1305), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1337), .B(new_n1292), .ZN(G402));
endmodule


