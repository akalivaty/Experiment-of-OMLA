

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;

  XNOR2_X1 U325 ( .A(n421), .B(n420), .ZN(n422) );
  NOR2_X1 U326 ( .A1(n410), .A2(n409), .ZN(n521) );
  XNOR2_X1 U327 ( .A(n415), .B(KEYINPUT37), .ZN(n416) );
  XNOR2_X1 U328 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U329 ( .A(n315), .B(n314), .Z(n522) );
  XOR2_X1 U330 ( .A(G211GAT), .B(KEYINPUT21), .Z(n293) );
  OR2_X1 U331 ( .A1(n556), .A2(n555), .ZN(n294) );
  INV_X1 U332 ( .A(KEYINPUT85), .ZN(n373) );
  XNOR2_X1 U333 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U334 ( .A(n374), .B(n373), .ZN(n375) );
  INV_X1 U335 ( .A(n423), .ZN(n426) );
  XNOR2_X1 U336 ( .A(n376), .B(n375), .ZN(n380) );
  NOR2_X1 U337 ( .A1(n562), .A2(n561), .ZN(n579) );
  INV_X1 U338 ( .A(KEYINPUT98), .ZN(n415) );
  XNOR2_X1 U339 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U340 ( .A(n417), .B(n416), .ZN(n496) );
  NOR2_X1 U341 ( .A1(n567), .A2(n566), .ZN(n576) );
  XOR2_X1 U342 ( .A(n450), .B(KEYINPUT38), .Z(n480) );
  XNOR2_X1 U343 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U344 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n296) );
  XNOR2_X1 U346 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U348 ( .A(KEYINPUT19), .B(n297), .ZN(n366) );
  INV_X1 U349 ( .A(n366), .ZN(n315) );
  XOR2_X1 U350 ( .A(KEYINPUT65), .B(KEYINPUT82), .Z(n299) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U353 ( .A(G176GAT), .B(G190GAT), .Z(n301) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G15GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n313) );
  XOR2_X1 U357 ( .A(G120GAT), .B(G71GAT), .Z(n430) );
  XOR2_X1 U358 ( .A(n430), .B(KEYINPUT20), .Z(n305) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U361 ( .A(n306), .B(G99GAT), .Z(n311) );
  XOR2_X1 U362 ( .A(KEYINPUT80), .B(G134GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(KEYINPUT81), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(KEYINPUT0), .B(n309), .Z(n392) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(n392), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n317) );
  XNOR2_X1 U370 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(G36GAT), .B(G190GAT), .Z(n363) );
  XOR2_X1 U373 ( .A(n318), .B(n363), .Z(n320) );
  XNOR2_X1 U374 ( .A(G134GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n330) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n368) );
  INV_X1 U377 ( .A(G85GAT), .ZN(n321) );
  NAND2_X1 U378 ( .A1(KEYINPUT72), .A2(n321), .ZN(n324) );
  INV_X1 U379 ( .A(KEYINPUT72), .ZN(n322) );
  NAND2_X1 U380 ( .A1(n322), .A2(G85GAT), .ZN(n323) );
  NAND2_X1 U381 ( .A1(n324), .A2(n323), .ZN(n326) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n421) );
  XOR2_X1 U384 ( .A(n368), .B(n421), .Z(n328) );
  NAND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U387 ( .A(n330), .B(n329), .Z(n338) );
  XOR2_X1 U388 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n332) );
  XNOR2_X1 U389 ( .A(G43GAT), .B(G29GAT), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U391 ( .A(KEYINPUT8), .B(n333), .Z(n445) );
  XOR2_X1 U392 ( .A(KEYINPUT66), .B(KEYINPUT75), .Z(n335) );
  XNOR2_X1 U393 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n445), .B(n336), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n549) );
  XNOR2_X1 U397 ( .A(n549), .B(KEYINPUT36), .ZN(n595) );
  XOR2_X1 U398 ( .A(G211GAT), .B(G155GAT), .Z(n340) );
  XNOR2_X1 U399 ( .A(G183GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U401 ( .A(n341), .B(G127GAT), .Z(n343) );
  XOR2_X1 U402 ( .A(G15GAT), .B(KEYINPUT70), .Z(n435) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(n435), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n356) );
  XOR2_X1 U405 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n345) );
  NAND2_X1 U406 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(G57GAT), .B(KEYINPUT13), .Z(n424) );
  XOR2_X1 U409 ( .A(n346), .B(n424), .Z(n354) );
  XOR2_X1 U410 ( .A(G64GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(G8GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n350) );
  XNOR2_X1 U414 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n591) );
  INV_X1 U419 ( .A(n591), .ZN(n545) );
  XNOR2_X1 U420 ( .A(G197GAT), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n293), .B(n357), .ZN(n369) );
  XOR2_X1 U422 ( .A(KEYINPUT88), .B(n369), .Z(n359) );
  NAND2_X1 U423 ( .A1(G226GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n362) );
  XOR2_X1 U425 ( .A(G64GAT), .B(G92GAT), .Z(n361) );
  XNOR2_X1 U426 ( .A(G176GAT), .B(G204GAT), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n423) );
  XOR2_X1 U428 ( .A(n362), .B(n423), .Z(n365) );
  XOR2_X1 U429 ( .A(G169GAT), .B(G8GAT), .Z(n436) );
  XNOR2_X1 U430 ( .A(n436), .B(n363), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U432 ( .A(n367), .B(n366), .Z(n476) );
  NAND2_X1 U433 ( .A1(n476), .A2(n522), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n371) );
  AND2_X1 U435 ( .A1(G228GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n376) );
  XNOR2_X1 U437 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n372), .B(KEYINPUT2), .ZN(n388) );
  XNOR2_X1 U439 ( .A(n388), .B(KEYINPUT23), .ZN(n374) );
  XOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n378) );
  XNOR2_X1 U441 ( .A(G106GAT), .B(G204GAT), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U443 ( .A(n380), .B(n379), .Z(n382) );
  XOR2_X1 U444 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XOR2_X1 U445 ( .A(G148GAT), .B(G78GAT), .Z(n429) );
  XNOR2_X1 U446 ( .A(n438), .B(n429), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n563) );
  NAND2_X1 U448 ( .A1(n383), .A2(n563), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n384), .B(KEYINPUT89), .ZN(n385) );
  XNOR2_X1 U450 ( .A(KEYINPUT25), .B(n385), .ZN(n387) );
  INV_X1 U451 ( .A(n476), .ZN(n552) );
  XOR2_X1 U452 ( .A(n552), .B(KEYINPUT27), .Z(n407) );
  NOR2_X1 U453 ( .A1(n563), .A2(n522), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n386), .B(KEYINPUT26), .ZN(n580) );
  NAND2_X1 U455 ( .A1(n407), .A2(n580), .ZN(n534) );
  NAND2_X1 U456 ( .A1(n387), .A2(n534), .ZN(n406) );
  XOR2_X1 U457 ( .A(G162GAT), .B(n388), .Z(n390) );
  XOR2_X1 U458 ( .A(G113GAT), .B(G1GAT), .Z(n437) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(n437), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n392), .B(n391), .ZN(n405) );
  XOR2_X1 U462 ( .A(G85GAT), .B(G148GAT), .Z(n394) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(G120GAT), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U465 ( .A(KEYINPUT86), .B(G57GAT), .Z(n396) );
  XNOR2_X1 U466 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n395) );
  XNOR2_X1 U467 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U468 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U469 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n400) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U472 ( .A(KEYINPUT1), .B(n401), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n562) );
  INV_X1 U475 ( .A(n562), .ZN(n497) );
  NAND2_X1 U476 ( .A1(n406), .A2(n497), .ZN(n412) );
  INV_X1 U477 ( .A(n407), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n563), .B(KEYINPUT28), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n408), .B(KEYINPUT67), .ZN(n479) );
  INV_X1 U480 ( .A(n479), .ZN(n504) );
  NAND2_X1 U481 ( .A1(n562), .A2(n504), .ZN(n409) );
  INV_X1 U482 ( .A(n522), .ZN(n566) );
  NAND2_X1 U483 ( .A1(n521), .A2(n566), .ZN(n411) );
  NAND2_X1 U484 ( .A1(n412), .A2(n411), .ZN(n457) );
  NAND2_X1 U485 ( .A1(n545), .A2(n457), .ZN(n413) );
  XOR2_X1 U486 ( .A(KEYINPUT97), .B(n413), .Z(n414) );
  NOR2_X1 U487 ( .A1(n595), .A2(n414), .ZN(n417) );
  NAND2_X1 U488 ( .A1(G230GAT), .A2(G233GAT), .ZN(n419) );
  INV_X1 U489 ( .A(KEYINPUT32), .ZN(n418) );
  XOR2_X1 U490 ( .A(KEYINPUT31), .B(n422), .Z(n428) );
  XNOR2_X1 U491 ( .A(n424), .B(KEYINPUT33), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n587) );
  XOR2_X1 U494 ( .A(KEYINPUT68), .B(G197GAT), .Z(n434) );
  XNOR2_X1 U495 ( .A(G50GAT), .B(G36GAT), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U497 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n442) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U504 ( .A(n445), .B(KEYINPUT29), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U506 ( .A(n449), .B(n448), .Z(n583) );
  INV_X1 U507 ( .A(n583), .ZN(n536) );
  NOR2_X1 U508 ( .A1(n587), .A2(n536), .ZN(n460) );
  NAND2_X1 U509 ( .A1(n496), .A2(n460), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n522), .A2(n480), .ZN(n454) );
  XOR2_X1 U511 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n452) );
  XNOR2_X1 U512 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n591), .A2(n549), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT79), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(KEYINPUT16), .ZN(n458) );
  NAND2_X1 U516 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U517 ( .A(KEYINPUT90), .B(n459), .Z(n484) );
  NAND2_X1 U518 ( .A1(n460), .A2(n484), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT91), .B(n461), .ZN(n470) );
  NAND2_X1 U520 ( .A1(n470), .A2(n562), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT34), .ZN(n463) );
  XNOR2_X1 U522 ( .A(G1GAT), .B(n463), .ZN(G1324GAT) );
  NAND2_X1 U523 ( .A1(n476), .A2(n470), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n466) );
  XNOR2_X1 U526 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U528 ( .A(KEYINPUT92), .B(n467), .Z(n469) );
  NAND2_X1 U529 ( .A1(n470), .A2(n522), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(G1326GAT) );
  XOR2_X1 U531 ( .A(G22GAT), .B(KEYINPUT95), .Z(n472) );
  NAND2_X1 U532 ( .A1(n470), .A2(n479), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(G1327GAT) );
  NAND2_X1 U534 ( .A1(n562), .A2(n480), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U537 ( .A(G29GAT), .B(n475), .ZN(G1328GAT) );
  XOR2_X1 U538 ( .A(G36GAT), .B(KEYINPUT99), .Z(n478) );
  NAND2_X1 U539 ( .A1(n480), .A2(n476), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(G1329GAT) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT102), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G50GAT), .B(n482), .ZN(G1331GAT) );
  XNOR2_X1 U544 ( .A(KEYINPUT41), .B(n587), .ZN(n539) );
  NOR2_X1 U545 ( .A1(n539), .A2(n583), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n483), .B(KEYINPUT104), .ZN(n495) );
  NAND2_X1 U547 ( .A1(n495), .A2(n484), .ZN(n490) );
  NOR2_X1 U548 ( .A1(n497), .A2(n490), .ZN(n486) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n485) );
  XNOR2_X1 U550 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U551 ( .A(G57GAT), .B(n487), .ZN(G1332GAT) );
  NOR2_X1 U552 ( .A1(n552), .A2(n490), .ZN(n488) );
  XOR2_X1 U553 ( .A(G64GAT), .B(n488), .Z(G1333GAT) );
  NOR2_X1 U554 ( .A1(n566), .A2(n490), .ZN(n489) );
  XOR2_X1 U555 ( .A(G71GAT), .B(n489), .Z(G1334GAT) );
  NOR2_X1 U556 ( .A1(n490), .A2(n504), .ZN(n494) );
  XOR2_X1 U557 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n492) );
  XNOR2_X1 U558 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n491) );
  XNOR2_X1 U559 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U560 ( .A(n494), .B(n493), .ZN(G1335GAT) );
  NAND2_X1 U561 ( .A1(n496), .A2(n495), .ZN(n503) );
  NOR2_X1 U562 ( .A1(n497), .A2(n503), .ZN(n498) );
  XOR2_X1 U563 ( .A(G85GAT), .B(n498), .Z(G1336GAT) );
  NOR2_X1 U564 ( .A1(n552), .A2(n503), .ZN(n500) );
  XNOR2_X1 U565 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U567 ( .A(G92GAT), .B(n501), .ZN(G1337GAT) );
  NOR2_X1 U568 ( .A1(n566), .A2(n503), .ZN(n502) );
  XOR2_X1 U569 ( .A(G99GAT), .B(n502), .Z(G1338GAT) );
  NOR2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT44), .B(n505), .Z(n506) );
  XNOR2_X1 U572 ( .A(G106GAT), .B(n506), .ZN(G1339GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n511) );
  NOR2_X1 U574 ( .A1(n536), .A2(n539), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n507), .B(KEYINPUT46), .ZN(n508) );
  NOR2_X1 U576 ( .A1(n508), .A2(n591), .ZN(n509) );
  NAND2_X1 U577 ( .A1(n509), .A2(n549), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n518) );
  XOR2_X1 U579 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n513) );
  NOR2_X1 U580 ( .A1(n545), .A2(n595), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(n514) );
  NOR2_X1 U582 ( .A1(n587), .A2(n514), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(KEYINPUT111), .ZN(n516) );
  NOR2_X1 U584 ( .A1(n583), .A2(n516), .ZN(n517) );
  NOR2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U586 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n556) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U589 ( .A1(n556), .A2(n523), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n531), .A2(n583), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT112), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  INV_X1 U594 ( .A(n539), .ZN(n569) );
  NAND2_X1 U595 ( .A1(n531), .A2(n569), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n529) );
  NAND2_X1 U598 ( .A1(n531), .A2(n591), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n533) );
  INV_X1 U602 ( .A(n549), .ZN(n575) );
  NAND2_X1 U603 ( .A1(n531), .A2(n575), .ZN(n532) );
  XNOR2_X1 U604 ( .A(n533), .B(n532), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n556), .A2(n534), .ZN(n535) );
  NAND2_X1 U606 ( .A1(n562), .A2(n535), .ZN(n548) );
  NOR2_X1 U607 ( .A1(n536), .A2(n548), .ZN(n537) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(n537), .Z(n538) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n539), .A2(n548), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n541) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n540) );
  XNOR2_X1 U613 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U614 ( .A(KEYINPUT52), .B(n542), .ZN(n543) );
  XNOR2_X1 U615 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n545), .A2(n548), .ZN(n547) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n546) );
  XNOR2_X1 U618 ( .A(n547), .B(n546), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(n550), .Z(n551) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n551), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n565) );
  XOR2_X1 U623 ( .A(KEYINPUT119), .B(n552), .Z(n555) );
  INV_X1 U624 ( .A(KEYINPUT121), .ZN(n553) );
  OR2_X1 U625 ( .A1(n555), .A2(n553), .ZN(n554) );
  OR2_X1 U626 ( .A1(n556), .A2(n554), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n553), .A2(n294), .ZN(n557) );
  NAND2_X1 U628 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U629 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n559) );
  XNOR2_X1 U630 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n579), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n576), .A2(n583), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .Z(n571) );
  NAND2_X1 U636 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NAND2_X1 U640 ( .A1(n591), .A2(n576), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n585) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U647 ( .A(KEYINPUT124), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n594) );
  NAND2_X1 U649 ( .A1(n583), .A2(n594), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(n586), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n594), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U655 ( .A(G204GAT), .B(n590), .Z(G1353GAT) );
  NAND2_X1 U656 ( .A1(n594), .A2(n591), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(KEYINPUT126), .ZN(n593) );
  XNOR2_X1 U658 ( .A(G211GAT), .B(n593), .ZN(G1354GAT) );
  INV_X1 U659 ( .A(n594), .ZN(n596) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U661 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

