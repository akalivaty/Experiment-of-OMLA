//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  XOR2_X1   g0007(.A(KEYINPUT65), .B(G238), .Z(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n207), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n207), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n217), .B(new_n220), .C1(new_n223), .C2(new_n225), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(KEYINPUT17), .ZN(new_n244));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n221), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(KEYINPUT70), .A3(new_n221), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT71), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n222), .A2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT79), .ZN(new_n261));
  INV_X1    g0061(.A(new_n253), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n255), .A2(new_n261), .B1(new_n262), .B2(new_n256), .ZN(new_n263));
  XNOR2_X1  g0063(.A(G58), .B(G68), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n267), .B(G20), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT77), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n270), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT77), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n222), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n272), .B1(new_n278), .B2(new_n267), .ZN(new_n279));
  OAI211_X1 g0079(.A(KEYINPUT16), .B(new_n266), .C1(new_n279), .C2(new_n209), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n281));
  NOR2_X1   g0081(.A1(new_n274), .A2(new_n275), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n267), .B1(new_n282), .B2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n269), .A2(new_n271), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n209), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n266), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n281), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n250), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n280), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n263), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G33), .A3(G41), .ZN(new_n296));
  INV_X1    g0096(.A(new_n221), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n221), .B1(KEYINPUT68), .B2(new_n293), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(KEYINPUT69), .A3(new_n296), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n292), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G1), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G41), .B2(G45), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n300), .A2(new_n302), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G232), .A3(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G87), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT80), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n269), .A2(new_n271), .A3(G226), .A4(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n269), .A2(new_n271), .A3(G223), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n297), .A2(new_n293), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT81), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n307), .A2(new_n309), .A3(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n312), .A2(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n244), .B1(new_n291), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n325), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n322), .B(KEYINPUT81), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n329), .A2(G200), .B1(new_n330), .B2(new_n311), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(KEYINPUT17), .A3(new_n290), .A4(new_n263), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n307), .A2(new_n309), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(new_n324), .B1(new_n325), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n291), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n334), .B1(new_n291), .B2(new_n338), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT82), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n291), .A2(new_n338), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT18), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT82), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(new_n339), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n333), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n255), .A2(G50), .A3(new_n259), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(G150), .ZN(new_n350));
  INV_X1    g0150(.A(new_n265), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n222), .A2(G33), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n349), .B1(new_n350), .B2(new_n351), .C1(new_n256), .C2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n289), .B1(new_n201), .B2(new_n262), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n355), .B(KEYINPUT9), .Z(new_n356));
  INV_X1    g0156(.A(G226), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n308), .A2(new_n305), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n284), .A2(new_n317), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G223), .B1(G77), .B2(new_n284), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n284), .A2(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G222), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n307), .B1(new_n357), .B2(new_n358), .C1(new_n363), .C2(new_n320), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G200), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n364), .A2(new_n310), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(KEYINPUT74), .A3(G200), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n356), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT73), .A4(new_n369), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n372), .C1(new_n356), .C2(new_n370), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n364), .A2(G179), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n364), .A2(new_n337), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n355), .A3(new_n378), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n253), .A2(G68), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT12), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n209), .ZN(new_n383));
  INV_X1    g0183(.A(G77), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n352), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n289), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n259), .A2(G68), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n386), .A2(new_n387), .B1(new_n254), .B2(new_n388), .ZN(new_n389));
  AOI211_X1 g0189(.A(new_n382), .B(new_n389), .C1(new_n387), .C2(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n391), .B(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n361), .B2(G226), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n282), .A2(G232), .A3(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n321), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n308), .A2(G238), .A3(new_n305), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n307), .A3(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n390), .B1(new_n402), .B2(new_n310), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n326), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(G169), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n400), .A2(G179), .A3(new_n401), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT14), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n409), .A3(G169), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n390), .B(KEYINPUT76), .Z(new_n412));
  AOI21_X1  g0212(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n352), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n256), .A2(new_n351), .B1(new_n222), .B2(new_n384), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n289), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n259), .A2(G77), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n417), .B1(G77), .B2(new_n253), .C1(new_n254), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n282), .A2(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G107), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n420), .A2(new_n208), .B1(new_n421), .B2(new_n282), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n282), .A2(G232), .A3(new_n317), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n321), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G244), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n307), .C1(new_n425), .C2(new_n358), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n419), .B1(new_n426), .B2(G200), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n310), .B2(new_n426), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n337), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n419), .C1(G179), .C2(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g0231(.A(new_n431), .B(KEYINPUT72), .Z(new_n432));
  AND4_X1   g0232(.A1(new_n347), .A2(new_n380), .A3(new_n413), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n269), .A2(new_n271), .A3(new_n222), .A4(G68), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT19), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n222), .A2(G33), .A3(G97), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n435), .A2(KEYINPUT87), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(G20), .B1(new_n393), .B2(KEYINPUT19), .ZN(new_n439));
  NOR3_X1   g0239(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n438), .B1(KEYINPUT87), .B2(new_n435), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(new_n289), .B1(new_n262), .B2(new_n414), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n304), .A2(G45), .ZN(new_n443));
  MUX2_X1   g0243(.A(G274), .B(G250), .S(new_n443), .Z(new_n444));
  NAND2_X1  g0244(.A1(new_n308), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G116), .ZN(new_n446));
  OR2_X1    g0246(.A1(G238), .A2(G1698), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n425), .A2(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n449), .B2(new_n284), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n321), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G200), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n304), .A2(G33), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n250), .A2(new_n253), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G87), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n442), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT88), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT88), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n442), .A2(new_n460), .A3(new_n453), .A4(new_n457), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n445), .A2(G190), .A3(new_n451), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n441), .A2(new_n289), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n455), .A2(new_n414), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n262), .A2(new_n414), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n452), .A2(G169), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n445), .A2(G179), .A3(new_n451), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n468), .B2(new_n469), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n467), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n222), .C1(G33), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G20), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n246), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n252), .A2(G20), .A3(new_n479), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n484), .C1(new_n479), .C2(new_n455), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G179), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n317), .ZN(new_n488));
  INV_X1    g0288(.A(G303), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n282), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n321), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n443), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n300), .B2(new_n302), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G270), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n308), .A2(G274), .A3(new_n495), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT89), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n490), .A2(new_n499), .A3(new_n321), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n492), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n486), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n485), .A3(G169), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT21), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(new_n485), .A3(new_n505), .A4(G169), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n485), .B1(new_n501), .B2(G200), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n310), .B2(new_n501), .ZN(new_n509));
  INV_X1    g0309(.A(new_n495), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n308), .A2(G257), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n498), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n359), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n361), .A2(KEYINPUT85), .A3(KEYINPUT4), .A4(G244), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(new_n317), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(new_n514), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n512), .B1(new_n321), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G190), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n498), .A2(new_n511), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n321), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n421), .B1(new_n283), .B2(new_n285), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n421), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n477), .A2(new_n421), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n533), .B2(KEYINPUT6), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n527), .B2(new_n528), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n289), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n455), .A2(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n253), .A2(new_n477), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT84), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n522), .A2(new_n526), .A3(new_n537), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n537), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n521), .A2(new_n335), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n525), .A2(new_n337), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n507), .A2(new_n509), .A3(new_n545), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT69), .B1(new_n301), .B2(new_n296), .ZN(new_n551));
  AND4_X1   g0351(.A1(KEYINPUT69), .A2(new_n294), .A3(new_n296), .A4(new_n297), .ZN(new_n552));
  OAI211_X1 g0352(.A(G264), .B(new_n510), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT91), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n496), .A2(new_n555), .A3(G264), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(new_n317), .ZN(new_n559));
  INV_X1    g0359(.A(G294), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n559), .C1(new_n268), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n321), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT92), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT92), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n561), .A2(new_n321), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n554), .C2(new_n556), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n498), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n498), .A2(new_n553), .A3(new_n562), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT90), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n568), .B(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n567), .A2(new_n326), .B1(new_n310), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n282), .A2(new_n222), .A3(G87), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT22), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n222), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n421), .A2(KEYINPUT23), .A3(G20), .ZN(new_n576));
  INV_X1    g0376(.A(new_n446), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n222), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g0379(.A(new_n579), .B(KEYINPUT24), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n289), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n262), .A2(new_n421), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n582), .B(KEYINPUT25), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n455), .A2(new_n421), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n571), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n585), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n580), .B2(new_n289), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n568), .B(KEYINPUT90), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n555), .B1(new_n496), .B2(G264), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n562), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n564), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n557), .A2(KEYINPUT92), .A3(new_n562), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(G179), .A3(new_n498), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n589), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT93), .B1(new_n587), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n591), .B1(new_n567), .B2(new_n335), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n586), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT93), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n603), .C1(new_n586), .C2(new_n571), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR4_X1   g0405(.A1(new_n434), .A2(new_n475), .A3(new_n550), .A4(new_n605), .ZN(G372));
  NOR2_X1   g0406(.A1(new_n340), .A2(new_n341), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n410), .A2(new_n408), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n409), .B1(new_n402), .B2(G169), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n412), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n405), .B2(new_n430), .ZN(new_n612));
  INV_X1    g0412(.A(new_n333), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n375), .A2(new_n376), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n379), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n467), .A2(new_n470), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n442), .A2(new_n453), .A3(new_n457), .A4(new_n462), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n549), .A2(new_n620), .A3(KEYINPUT26), .ZN(new_n621));
  INV_X1    g0421(.A(new_n549), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n463), .A3(new_n474), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n623), .B2(KEYINPUT26), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n545), .A2(new_n549), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n619), .C1(new_n586), .C2(new_n571), .ZN(new_n626));
  INV_X1    g0426(.A(new_n507), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n599), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n618), .B(new_n624), .C1(new_n626), .C2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n617), .B1(new_n434), .B2(new_n630), .ZN(G369));
  INV_X1    g0431(.A(new_n252), .ZN(new_n632));
  OR3_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .A3(G20), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT27), .B1(new_n632), .B2(G20), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n485), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n507), .A2(new_n509), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n507), .B2(new_n638), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  INV_X1    g0441(.A(new_n637), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n600), .B(new_n604), .C1(new_n589), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n599), .A2(new_n637), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n507), .A2(new_n637), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n600), .A2(new_n604), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n599), .A2(new_n642), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n645), .A2(new_n649), .ZN(G399));
  INV_X1    g0450(.A(new_n218), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G41), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n440), .A2(new_n479), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(G1), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n653), .A2(new_n224), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(KEYINPUT94), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(KEYINPUT94), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT29), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n629), .A2(new_n661), .A3(new_n642), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n545), .A2(new_n549), .A3(new_n619), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n587), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n602), .A2(new_n507), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n467), .B2(new_n470), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n549), .A2(new_n620), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(KEYINPUT26), .B2(new_n623), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n637), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n662), .B1(new_n671), .B2(new_n661), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n445), .A2(G179), .A3(new_n451), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n490), .A2(new_n499), .A3(new_n321), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n499), .B1(new_n490), .B2(new_n321), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(G270), .A2(new_n496), .B1(new_n303), .B2(new_n495), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n525), .ZN(new_n679));
  AOI211_X1 g0479(.A(KEYINPUT96), .B(KEYINPUT30), .C1(new_n597), .C2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT96), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n501), .A2(new_n469), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n521), .B(new_n682), .C1(new_n563), .C2(new_n566), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT97), .ZN(new_n687));
  INV_X1    g0487(.A(new_n567), .ZN(new_n688));
  AOI21_X1  g0488(.A(G179), .B1(new_n445), .B2(new_n451), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n501), .A2(KEYINPUT95), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT95), .B1(new_n501), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n525), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n688), .A2(new_n693), .B1(new_n684), .B2(new_n683), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n686), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n563), .A2(new_n566), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n682), .A2(new_n521), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n684), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT96), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n683), .A2(new_n681), .A3(new_n684), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n683), .ZN(new_n702));
  INV_X1    g0502(.A(new_n692), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n521), .B1(new_n703), .B2(new_n690), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n702), .A2(KEYINPUT30), .B1(new_n704), .B2(new_n567), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT97), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n637), .B1(new_n695), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n698), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n642), .A2(new_n708), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n550), .A2(new_n475), .A3(new_n637), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n600), .A2(new_n713), .A3(new_n604), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n672), .B1(G330), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n660), .B1(new_n716), .B2(G1), .ZN(G364));
  INV_X1    g0517(.A(new_n641), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n251), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n304), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n652), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n640), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n218), .A2(new_n282), .ZN(new_n725));
  INV_X1    g0525(.A(G355), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n726), .B1(G116), .B2(new_n218), .ZN(new_n727));
  INV_X1    g0527(.A(G45), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n239), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n276), .A2(new_n277), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n218), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n728), .B2(new_n225), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n727), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n221), .B1(G20), .B2(new_n337), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n722), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n222), .A2(new_n326), .A3(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n310), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n421), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(G87), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n222), .A2(new_n335), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n310), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n748), .B1(new_n201), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n750), .A2(G190), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n744), .B(new_n753), .C1(G68), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G20), .A3(new_n335), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G159), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT32), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n335), .A2(new_n326), .A3(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n759), .A2(KEYINPUT32), .B1(G97), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n749), .A2(G190), .A3(new_n326), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n282), .B1(new_n764), .B2(new_n202), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n749), .A2(new_n756), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G77), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n755), .A2(new_n760), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G317), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT33), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(KEYINPUT33), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n754), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n762), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n773), .B1(new_n560), .B2(new_n774), .C1(new_n489), .C2(new_n745), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n282), .B1(G329), .B2(new_n758), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n776), .B1(new_n777), .B2(new_n766), .C1(new_n778), .C2(new_n764), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n751), .A2(G326), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n743), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n775), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n741), .B1(new_n785), .B2(new_n738), .ZN(new_n786));
  INV_X1    g0586(.A(new_n737), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n640), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n724), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  NAND2_X1  g0590(.A1(new_n715), .A2(G330), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n419), .A2(new_n637), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n428), .A2(new_n430), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT99), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n430), .A2(new_n642), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n630), .B2(new_n637), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n629), .A2(new_n642), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n722), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n791), .B2(new_n801), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n738), .A2(new_n735), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n722), .B1(G77), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n754), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n781), .A2(new_n807), .B1(new_n752), .B2(new_n489), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G107), .B2(new_n746), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n762), .A2(G97), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n764), .A2(new_n560), .B1(new_n757), .B2(new_n777), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n282), .B(new_n811), .C1(G116), .C2(new_n767), .ZN(new_n812));
  INV_X1    g0612(.A(new_n743), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G87), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n809), .A2(new_n810), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n764), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G143), .B1(new_n767), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n752), .B2(new_n818), .C1(new_n350), .C2(new_n807), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n731), .B1(G132), .B2(new_n758), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n743), .A2(new_n209), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n202), .B2(new_n774), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G50), .B2(new_n746), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n819), .A2(new_n820), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n815), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n806), .B1(new_n829), .B2(new_n738), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n794), .B(new_n795), .C1(new_n430), .C2(new_n642), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n736), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n803), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G384));
  NOR2_X1   g0634(.A1(new_n719), .A2(new_n304), .ZN(new_n835));
  INV_X1    g0635(.A(new_n405), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n412), .A2(new_n637), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n611), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n412), .B(new_n637), .C1(new_n411), .C2(new_n405), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n798), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT40), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n331), .A2(new_n290), .A3(new_n263), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n255), .A2(new_n261), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n262), .A2(new_n256), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n266), .B1(new_n279), .B2(new_n209), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT100), .B(new_n266), .C1(new_n279), .C2(new_n209), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n281), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n280), .A2(new_n289), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n845), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n338), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n635), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n635), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n291), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n842), .A2(new_n343), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n855), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n861), .B(KEYINPUT38), .C1(new_n347), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n842), .A2(new_n343), .A3(new_n858), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(new_n859), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n858), .B1(new_n613), .B2(new_n607), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n841), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n711), .B1(new_n695), .B2(new_n706), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n714), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n687), .B1(new_n686), .B2(new_n694), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n701), .A2(KEYINPUT97), .A3(new_n705), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT31), .B1(new_n874), .B2(new_n637), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n840), .B(new_n869), .C1(new_n871), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n642), .B1(new_n872), .B2(new_n873), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n870), .B(new_n714), .C1(new_n878), .C2(KEYINPUT31), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n840), .A4(new_n869), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n861), .B1(new_n347), .B2(new_n862), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n864), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n863), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n879), .A2(new_n884), .A3(new_n840), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n877), .A2(new_n881), .B1(new_n841), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n433), .A2(new_n879), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  INV_X1    g0689(.A(G330), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n838), .A2(new_n839), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n430), .A2(new_n637), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n800), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n897), .A2(new_n884), .B1(new_n608), .B2(new_n635), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n863), .A2(new_n868), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n411), .A2(new_n412), .A3(new_n642), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n901), .B(new_n903), .C1(new_n884), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n616), .B1(new_n672), .B2(new_n433), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n905), .B(new_n906), .Z(new_n907));
  AOI21_X1  g0707(.A(new_n835), .B1(new_n892), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n892), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n910), .A2(G116), .A3(new_n223), .A4(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  OAI21_X1  g0713(.A(G77), .B1(new_n202), .B2(new_n209), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n914), .A2(new_n224), .B1(G50), .B2(new_n209), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(G1), .A3(new_n251), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT102), .Z(G367));
  NAND2_X1  g0718(.A1(new_n442), .A2(new_n457), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n637), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n618), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT103), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n618), .A3(new_n619), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n546), .A2(new_n637), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n625), .A2(new_n926), .B1(new_n622), .B2(new_n637), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n647), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n625), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n549), .B1(new_n929), .B2(new_n602), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n928), .A2(KEYINPUT42), .B1(new_n642), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n925), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n935), .ZN(new_n939));
  INV_X1    g0739(.A(new_n933), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n940), .A2(new_n931), .B1(KEYINPUT43), .B2(new_n924), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n937), .A2(new_n935), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n645), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n927), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n938), .A2(new_n943), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n944), .B2(new_n927), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n652), .B(KEYINPUT41), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n649), .A2(new_n927), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n649), .A2(new_n927), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT44), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n645), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n951), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n950), .B(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT44), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n953), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n944), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n646), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n643), .A2(new_n644), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n647), .B1(new_n962), .B2(KEYINPUT107), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n718), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n967), .A2(new_n641), .A3(new_n647), .A4(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n955), .A2(new_n960), .A3(new_n969), .A4(new_n716), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n949), .B1(new_n970), .B2(new_n716), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n946), .B(new_n948), .C1(new_n971), .C2(new_n721), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n739), .B1(new_n218), .B2(new_n414), .C1(new_n732), .C2(new_n234), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n722), .ZN(new_n974));
  INV_X1    g0774(.A(new_n738), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n743), .A2(new_n384), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n284), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT109), .Z(new_n978));
  OAI22_X1  g0778(.A1(new_n766), .A2(new_n201), .B1(new_n757), .B2(new_n818), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G150), .B2(new_n816), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G143), .A2(new_n751), .B1(new_n754), .B2(G159), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n746), .A2(G58), .B1(new_n762), .B2(G68), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT108), .B(G311), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n560), .A2(new_n807), .B1(new_n752), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G97), .B2(new_n813), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n764), .A2(new_n489), .B1(new_n766), .B2(new_n781), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G317), .B2(new_n758), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n730), .B1(G107), .B2(new_n762), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n746), .A2(G116), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n986), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  OAI221_X1 g0794(.A(new_n974), .B1(new_n975), .B2(new_n994), .C1(new_n924), .C2(new_n787), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n972), .A2(new_n996), .ZN(G387));
  OR2_X1    g0797(.A1(new_n969), .A2(new_n716), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n653), .B1(new_n969), .B2(new_n716), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n643), .A2(new_n644), .A3(new_n737), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n231), .A2(G45), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1001), .A2(new_n732), .B1(new_n655), .B2(new_n725), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n256), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT50), .B1(new_n256), .B2(G50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n655), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1002), .A2(new_n1006), .B1(new_n421), .B2(new_n651), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n722), .B1(new_n1007), .B2(new_n740), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n816), .A2(G317), .B1(new_n767), .B2(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n752), .B2(new_n778), .C1(new_n807), .C2(new_n984), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n746), .A2(G294), .B1(new_n762), .B2(G283), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n743), .A2(new_n479), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n730), .B(new_n1019), .C1(G326), .C2(new_n758), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n754), .A2(new_n257), .B1(new_n767), .B2(G68), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT112), .Z(new_n1023));
  INV_X1    g0823(.A(G159), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n752), .A2(new_n1024), .B1(new_n477), .B2(new_n743), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n774), .A2(new_n414), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n745), .A2(new_n384), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n816), .A2(G50), .B1(G150), .B2(new_n758), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n730), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1021), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1008), .B1(new_n1031), .B2(new_n738), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n998), .A2(new_n999), .B1(new_n1000), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n720), .B1(new_n966), .B2(new_n968), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(G393));
  NAND3_X1  g0836(.A1(new_n955), .A2(new_n721), .A3(new_n960), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n927), .A2(new_n737), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n739), .B1(new_n477), .B2(new_n218), .C1(new_n732), .C2(new_n242), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n722), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT113), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n774), .A2(new_n384), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n814), .B1(new_n209), .B2(new_n745), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G50), .C2(new_n754), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n752), .A2(new_n350), .B1(new_n1024), .B2(new_n764), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n767), .A2(new_n257), .B1(new_n758), .B2(G143), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n730), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n752), .A2(new_n770), .B1(new_n777), .B2(new_n764), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n754), .A2(G303), .B1(G116), .B2(new_n762), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n284), .B1(new_n757), .B2(new_n778), .C1(new_n766), .C2(new_n560), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n744), .B(new_n1054), .C1(G283), .C2(new_n746), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1038), .B(new_n1041), .C1(new_n975), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n970), .A2(new_n652), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n955), .A2(new_n960), .B1(new_n969), .B2(new_n716), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1037), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(G390));
  NAND2_X1  g0861(.A1(new_n714), .A2(new_n712), .ZN(new_n1062));
  OAI211_X1 g0862(.A(G330), .B(new_n831), .C1(new_n875), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n894), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n879), .A2(G330), .A3(new_n840), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n800), .A2(new_n896), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT115), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT115), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1067), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n711), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n872), .B2(new_n873), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n600), .A2(new_n604), .A3(new_n713), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n890), .B1(new_n1075), .B2(new_n709), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n893), .B1(new_n1076), .B2(new_n831), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n895), .B1(new_n671), .B2(new_n796), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1063), .B2(new_n894), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1068), .A2(new_n1071), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(new_n433), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n906), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1063), .A2(new_n894), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n901), .B1(new_n884), .B2(new_n900), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n903), .B2(new_n897), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n902), .B(new_n899), .C1(new_n1078), .C2(new_n894), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n1065), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n653), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1065), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1089), .B2(new_n1084), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1080), .A2(new_n1093), .A3(new_n1082), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n721), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n722), .B1(new_n257), .B2(new_n805), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n807), .A2(new_n818), .B1(new_n1024), .B2(new_n774), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G128), .B2(new_n751), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n745), .A2(new_n350), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n764), .A2(new_n1102), .B1(new_n757), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n767), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1099), .A2(new_n1101), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n282), .B1(new_n743), .B2(new_n201), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT116), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n764), .A2(new_n479), .B1(new_n757), .B2(new_n560), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n282), .B(new_n1111), .C1(G97), .C2(new_n767), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n748), .A3(new_n824), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1042), .B1(G283), .B2(new_n751), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n421), .B2(new_n807), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1108), .A2(new_n1110), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1097), .B1(new_n1116), .B2(new_n738), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1085), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n736), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1096), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1095), .A2(new_n1121), .ZN(G378));
  INV_X1    g0922(.A(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n355), .A2(new_n857), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n380), .B(new_n1124), .Z(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1126));
  XNOR2_X1  g0926(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n885), .A2(new_n841), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n893), .A2(new_n831), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1075), .B2(new_n709), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n880), .B1(new_n1131), .B2(new_n869), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n881), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n1129), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n905), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n905), .B1(new_n886), .B2(G330), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1128), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n886), .A2(G330), .A3(new_n905), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1127), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n720), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1128), .A2(new_n736), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1103), .A2(new_n752), .B1(new_n807), .B2(new_n1102), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n816), .A2(G128), .B1(new_n767), .B2(G137), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n745), .B2(new_n1105), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G150), .C2(new_n762), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(KEYINPUT59), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n813), .A2(G159), .ZN(new_n1151));
  AOI211_X1 g0951(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n764), .A2(new_n421), .B1(new_n766), .B2(new_n414), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n730), .A2(G41), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G283), .C2(new_n758), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n743), .A2(new_n202), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT117), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1027), .B1(G68), .B2(new_n762), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G97), .A2(new_n754), .B1(new_n751), .B2(G116), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT58), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1156), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1166));
  AND4_X1   g0966(.A1(new_n1153), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n722), .B1(G50), .B2(new_n805), .C1(new_n1167), .C2(new_n975), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1143), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1123), .B1(new_n1142), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1139), .A2(new_n1127), .A3(new_n1140), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1127), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n721), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1169), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(KEYINPUT118), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n840), .A2(new_n1076), .B1(new_n1063), .B2(new_n894), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1069), .B1(new_n1178), .B2(new_n1070), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1066), .A2(KEYINPUT115), .A3(new_n1067), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1082), .B1(new_n1181), .B2(new_n1090), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(KEYINPUT57), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1094), .A2(new_n1082), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n652), .C1(new_n1184), .C2(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1176), .A2(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n894), .A2(new_n735), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n722), .B1(G68), .B2(new_n805), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT119), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n807), .A2(new_n1105), .B1(new_n1024), .B2(new_n745), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G132), .B2(new_n751), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n816), .A2(G137), .B1(G128), .B2(new_n758), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n730), .A2(new_n1191), .A3(new_n1159), .A4(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n774), .A2(new_n201), .B1(new_n350), .B2(new_n766), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT121), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n745), .A2(new_n477), .B1(new_n489), .B2(new_n757), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT120), .Z(new_n1197));
  OAI22_X1  g0997(.A1(new_n479), .A2(new_n807), .B1(new_n752), .B2(new_n560), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n284), .B1(new_n766), .B2(new_n421), .C1(new_n781), .C2(new_n764), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1198), .A2(new_n976), .A3(new_n1026), .A4(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1193), .A2(new_n1195), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1189), .B1(new_n1201), .B2(new_n975), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT122), .Z(new_n1203));
  AOI22_X1  g1003(.A1(new_n1080), .A2(new_n721), .B1(new_n1187), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n949), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1083), .A2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1082), .B(new_n1177), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(G381));
  OR2_X1    g1008(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  INV_X1    g1011(.A(G390), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n833), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(G378), .A2(new_n1213), .A3(G387), .A4(G381), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1214), .ZN(G407));
  NAND2_X1  g1015(.A1(new_n636), .A2(G213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G378), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1209), .A2(new_n1210), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G407), .A2(new_n1218), .A3(G213), .ZN(G409));
  NAND3_X1  g1019(.A1(new_n1176), .A2(new_n1185), .A3(G378), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1120), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1184), .A2(new_n1205), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1207), .B1(new_n1083), .B2(KEYINPUT60), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1082), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n652), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1204), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1230), .A2(new_n833), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G384), .B(new_n1204), .C1(new_n1226), .C2(new_n1229), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1225), .A2(new_n1216), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT62), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1225), .A2(new_n1216), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1230), .A2(new_n833), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1238), .A2(new_n1232), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1238), .B2(new_n1232), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1225), .A2(new_n1245), .A3(new_n1234), .A4(new_n1216), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1236), .A2(new_n1243), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(G396), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n972), .A2(new_n996), .A3(G390), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G390), .B1(new_n972), .B2(new_n996), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1212), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n789), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1211), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n972), .A2(new_n996), .A3(G390), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1251), .A2(new_n1256), .A3(KEYINPUT125), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT125), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1254), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1251), .A2(new_n1256), .A3(KEYINPUT125), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1260), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1247), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1235), .A2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1225), .A2(KEYINPUT63), .A3(new_n1234), .A4(new_n1216), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(G405));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1234), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT127), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1220), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1176), .B2(new_n1185), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1277), .B(new_n1278), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1276), .A3(new_n1234), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1265), .A4(new_n1264), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(G402));
endmodule


