//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(new_n459));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n453), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n478), .B(new_n481), .C1(G136), .C2(new_n472), .ZN(G162));
  NAND2_X1  g057(.A1(new_n472), .A2(G138), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n472), .A2(new_n485), .A3(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT71), .B1(new_n489), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n490), .A2(new_n493), .A3(G2104), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  OAI21_X1  g092(.A(KEYINPUT72), .B1(new_n509), .B2(new_n508), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n502), .A2(new_n519), .A3(new_n503), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n524), .B1(new_n525), .B2(new_n514), .C1(new_n526), .C2(new_n512), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G168));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n520), .A3(G64), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n506), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n512), .A2(new_n532), .B1(new_n514), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n512), .A2(new_n536), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n518), .A2(new_n520), .A3(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n538), .B1(new_n541), .B2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n506), .B1(new_n539), .B2(new_n540), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n538), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  XNOR2_X1  g127(.A(KEYINPUT75), .B(G65), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n504), .A2(new_n553), .B1(G78), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n506), .ZN(new_n555));
  INV_X1    g130(.A(new_n512), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n514), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n514), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n518), .A2(new_n520), .ZN(new_n569));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n506), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  INV_X1    g147(.A(G49), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n512), .A2(new_n572), .B1(new_n514), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n506), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n512), .A2(new_n579), .B1(new_n514), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n521), .A2(G60), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n506), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT76), .B(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n512), .A2(new_n587), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n556), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n504), .A2(G66), .ZN(new_n596));
  INV_X1    g171(.A(G79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n501), .ZN(new_n598));
  INV_X1    g173(.A(new_n514), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n598), .A2(G651), .B1(new_n599), .B2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n564), .ZN(G297));
  XOR2_X1   g181(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n602), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n468), .A2(new_n473), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G2100), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT79), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n480), .A2(G123), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n472), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n489), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G2096), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(G2100), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n620), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT80), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(KEYINPUT17), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT81), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n655), .A2(new_n648), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n649), .A2(new_n648), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n654), .B(new_n657), .C1(new_n652), .C2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n663), .A2(new_n666), .A3(new_n670), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  XOR2_X1   g256(.A(KEYINPUT84), .B(G29), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(G25), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n480), .A2(G119), .ZN(new_n685));
  NOR2_X1   g260(.A1(G95), .A2(G2105), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT85), .Z(new_n687));
  INV_X1    g262(.A(G107), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n465), .B1(new_n688), .B2(G2105), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n687), .A2(new_n689), .B1(G131), .B2(new_n472), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n684), .B1(new_n692), .B2(new_n683), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT35), .B(G1991), .Z(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n575), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n696), .B2(G23), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT88), .B(G1971), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n698), .A2(new_n700), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n696), .A2(G6), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n582), .B2(new_n696), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n701), .A2(new_n705), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n695), .B1(KEYINPUT34), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n696), .A2(G24), .ZN(new_n713));
  NOR2_X1   g288(.A1(G290), .A2(KEYINPUT86), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n715));
  OAI21_X1  g290(.A(G16), .B1(new_n590), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n712), .B(new_n719), .C1(KEYINPUT34), .C2(new_n711), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n682), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G128), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(G116), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G2105), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G140), .B2(new_n472), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n729), .A2(KEYINPUT92), .A3(G29), .ZN(new_n730));
  AOI21_X1  g305(.A(KEYINPUT92), .B1(new_n729), .B2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n723), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT93), .B(G2067), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n547), .A2(new_n696), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n696), .B2(G19), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT91), .B(G1341), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n683), .A2(G35), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n683), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT29), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G2090), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(G2090), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n696), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n696), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT94), .Z(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n744), .A2(new_n745), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n480), .A2(G129), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n472), .A2(G141), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT26), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n473), .A2(G105), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n753), .A2(new_n754), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  MUX2_X1   g333(.A(G32), .B(new_n758), .S(G29), .Z(new_n759));
  XOR2_X1   g334(.A(KEYINPUT27), .B(G1996), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT24), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G34), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(G34), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n683), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G160), .B2(G29), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n766), .B1(new_n771), .B2(G2084), .C1(new_n625), .C2(new_n682), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n761), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n489), .A2(G103), .A3(G2104), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT25), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n468), .A2(G127), .ZN(new_n776));
  NAND2_X1  g351(.A1(G115), .A2(G2104), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n489), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n775), .B(new_n778), .C1(G139), .C2(new_n472), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G29), .B2(G33), .ZN(new_n781));
  INV_X1    g356(.A(G2072), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n781), .A2(new_n782), .B1(G2084), .B2(new_n771), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n773), .B(new_n783), .C1(new_n782), .C2(new_n781), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n696), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n696), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n696), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(G1961), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n683), .A2(G27), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n683), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G2078), .Z(new_n795));
  NAND4_X1  g370(.A1(new_n788), .A2(new_n791), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n602), .A2(new_n696), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G4), .B2(new_n696), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT89), .B(G1348), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT90), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n759), .A2(new_n760), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n798), .A2(new_n800), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n784), .A2(new_n796), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n721), .A2(new_n740), .A3(new_n752), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n512), .A2(new_n808), .B1(new_n514), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n518), .A2(new_n520), .A3(G67), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n810), .B1(new_n813), .B2(G651), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(G651), .ZN(new_n818));
  INV_X1    g393(.A(new_n810), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n543), .A2(new_n546), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n820), .A2(KEYINPUT95), .A3(new_n542), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n541), .A2(G651), .ZN(new_n824));
  INV_X1    g399(.A(new_n538), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(new_n826), .B2(new_n814), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n821), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT96), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(new_n821), .C1(new_n822), .C2(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n601), .A2(new_n608), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n815), .B1(new_n836), .B2(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n817), .B1(new_n837), .B2(new_n838), .ZN(G145));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n758), .B(new_n729), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n480), .A2(G130), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n472), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n489), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n841), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n691), .B(new_n616), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n496), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n488), .A2(new_n495), .A3(KEYINPUT97), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n487), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n779), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n850), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n625), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n840), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n860), .A2(KEYINPUT98), .A3(new_n864), .A4(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n862), .B2(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g446(.A(G868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n820), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n831), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT95), .B1(new_n820), .B2(new_n542), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n826), .A2(new_n823), .A3(new_n814), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n830), .B1(new_n877), .B2(new_n821), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n610), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n602), .A2(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n601), .A2(new_n564), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(new_n881), .B2(new_n882), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI22_X1  g462(.A1(new_n884), .A2(KEYINPUT99), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(KEYINPUT99), .B2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(G290), .A2(new_n582), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n590), .A2(G305), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n575), .B(G166), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n893), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n889), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n873), .B1(new_n900), .B2(new_n872), .ZN(G295));
  OAI21_X1  g476(.A(new_n873), .B1(new_n900), .B2(new_n872), .ZN(G331));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT103), .B1(new_n895), .B2(new_n896), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  INV_X1    g483(.A(new_n534), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n529), .A2(new_n530), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n506), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT101), .B1(new_n531), .B2(new_n534), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n911), .A2(G168), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G168), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n829), .A2(new_n831), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n832), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  AOI211_X1 g494(.A(new_n919), .B(new_n915), .C1(new_n829), .C2(new_n831), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n887), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n916), .A2(new_n883), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n917), .B1(new_n874), .B2(new_n878), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n907), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n919), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n832), .A2(KEYINPUT102), .A3(new_n917), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n887), .B1(new_n931), .B2(new_n916), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n926), .A2(new_n897), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n897), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n924), .B2(new_n925), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n929), .A2(new_n930), .B1(new_n879), .B2(new_n915), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n938), .B2(new_n887), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n916), .A2(new_n883), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n929), .B2(new_n930), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n887), .B1(new_n916), .B2(new_n925), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n906), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .A4(new_n928), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT104), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n923), .B2(new_n937), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n944), .A4(new_n943), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n935), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n927), .A2(new_n934), .A3(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n943), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n953), .B2(new_n955), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(G397));
  NAND3_X1  g534(.A1(new_n487), .A2(new_n853), .A3(new_n854), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT106), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n729), .A2(G2067), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n729), .A2(G2067), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n758), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n691), .B(new_n694), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(KEYINPUT107), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(KEYINPUT107), .B2(new_n973), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n590), .B(new_n718), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n601), .B(KEYINPUT121), .Z(new_n978));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n960), .A2(new_n980), .A3(new_n961), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n487), .B2(new_n497), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n981), .B(new_n963), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n963), .A2(new_n960), .A3(new_n961), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(G2067), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n983), .A2(new_n799), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT117), .B1(new_n984), .B2(G2067), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n979), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n799), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(new_n986), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n979), .A2(new_n990), .A3(new_n988), .A4(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT60), .B(new_n978), .C1(new_n989), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n988), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT118), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT60), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n987), .A2(new_n979), .A3(new_n988), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n601), .A2(KEYINPUT121), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n993), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n960), .A2(new_n961), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1004), .A2(KEYINPUT112), .B1(new_n980), .B2(new_n982), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n980), .B1(new_n960), .B2(new_n961), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT114), .B(G1956), .Z(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n498), .A2(new_n961), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n960), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n963), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1009), .A2(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n558), .B1(new_n1020), .B2(new_n562), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n563), .A2(KEYINPUT115), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n564), .A2(KEYINPUT57), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1028), .A3(new_n1024), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT119), .B1(new_n1019), .B2(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1010), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1032), .B(new_n1033), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1019), .A2(new_n1030), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1031), .A2(KEYINPUT61), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT61), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1036), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1030), .B1(new_n1042), .B2(new_n1034), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1015), .A2(new_n963), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n969), .A3(new_n1014), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n984), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1046), .A2(KEYINPUT120), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT120), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n547), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT59), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(new_n547), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1001), .A2(new_n1039), .A3(new_n1044), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n995), .A2(new_n602), .A3(new_n997), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1031), .A2(new_n1057), .A3(new_n1037), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1038), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1016), .B2(G2078), .ZN(new_n1062));
  INV_X1    g637(.A(G1961), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n983), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n962), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1045), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1068), .B2(KEYINPUT123), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(KEYINPUT123), .B2(new_n1068), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1002), .B1(new_n982), .B2(KEYINPUT45), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1062), .A2(new_n1072), .A3(new_n1064), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(KEYINPUT54), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT108), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n983), .B2(G2090), .ZN(new_n1077));
  INV_X1    g652(.A(G1971), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1016), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1002), .B1(new_n1012), .B2(KEYINPUT50), .ZN(new_n1080));
  INV_X1    g655(.A(G2090), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(KEYINPUT108), .A3(new_n1081), .A4(new_n981), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G166), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT55), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(G8), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n575), .A2(G1976), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n984), .A2(G8), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(KEYINPUT109), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n575), .A2(G1976), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n984), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(G1981), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n582), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT110), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n582), .A2(KEYINPUT110), .A3(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n578), .B1(new_n581), .B2(KEYINPUT111), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(KEYINPUT111), .B2(new_n581), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G1981), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1095), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(new_n1104), .A3(KEYINPUT49), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1107), .A2(new_n1108), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1087), .A2(new_n1094), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1005), .A2(new_n1081), .A3(new_n1008), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1084), .B1(new_n1111), .B2(new_n1079), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n1086), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n963), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1115), .B(new_n749), .C1(new_n1116), .C2(new_n962), .ZN(new_n1117));
  INV_X1    g692(.A(G2084), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1080), .A2(new_n1118), .A3(new_n981), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1115), .B1(new_n1121), .B2(new_n749), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G168), .A2(new_n1084), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(KEYINPUT51), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n749), .B1(new_n1116), .B2(new_n962), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT113), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(new_n1119), .A3(new_n1117), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1127), .B(G8), .C1(new_n1130), .C2(G286), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT122), .B(new_n1124), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT122), .B1(new_n1130), .B2(new_n1124), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1126), .B(new_n1131), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1073), .A2(G171), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1062), .A2(G301), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT54), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1075), .A2(new_n1114), .A3(new_n1135), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1138), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1143), .A2(KEYINPUT124), .A3(new_n1075), .A4(new_n1135), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1060), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1135), .A2(KEYINPUT62), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT125), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1135), .A2(KEYINPUT62), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1135), .A2(new_n1149), .A3(KEYINPUT62), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1109), .A2(new_n1094), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1152), .B(new_n1087), .C1(new_n1086), .C2(new_n1112), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(new_n1136), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G288), .A2(G1976), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1156), .A2(new_n1157), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1151), .A2(new_n1087), .B1(new_n1158), .B2(new_n1095), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1130), .A2(G8), .A3(G168), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1083), .A2(G8), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(new_n1086), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(new_n1160), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1164), .A2(new_n1087), .A3(new_n1152), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1159), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1155), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n977), .B1(new_n1145), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n975), .A2(new_n965), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n965), .A2(new_n718), .A3(new_n590), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT48), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1170), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n968), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n965), .B1(new_n1176), .B2(new_n758), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n965), .A2(new_n1178), .A3(new_n969), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1178), .B1(new_n965), .B2(new_n969), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT47), .Z(new_n1182));
  NAND2_X1  g757(.A1(new_n692), .A2(new_n694), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n966), .B1(new_n971), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1175), .B(new_n1182), .C1(new_n965), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1169), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g761(.A1(G227), .A2(new_n462), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n646), .A2(new_n680), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g765(.A1(new_n646), .A2(new_n680), .A3(KEYINPUT126), .A4(new_n1188), .ZN(new_n1192));
  AOI22_X1  g766(.A1(new_n868), .A2(new_n869), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n950), .A2(KEYINPUT127), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g768(.A(KEYINPUT127), .B1(new_n950), .B2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1195), .ZN(G308));
  NAND2_X1  g770(.A1(new_n950), .A2(new_n1193), .ZN(G225));
endmodule


