//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(G1gat), .ZN(new_n210));
  AOI21_X1  g009(.A(G8gat), .B1(new_n210), .B2(KEYINPUT94), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT16), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(G1gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n211), .B(new_n217), .Z(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(KEYINPUT15), .B(new_n219), .C1(new_n221), .C2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT92), .B1(new_n222), .B2(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(new_n221), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n219), .B(KEYINPUT15), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n218), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(KEYINPUT13), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n232), .B(KEYINPUT17), .ZN(new_n237));
  INV_X1    g036(.A(new_n218), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n232), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT95), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n236), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n244), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n208), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n239), .A2(new_n240), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n234), .A3(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n244), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n249), .A2(new_n207), .A3(new_n250), .A4(new_n236), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G141gat), .B(G148gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(KEYINPUT2), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT80), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(G155gat), .A3(G162gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G155gat), .ZN(new_n261));
  INV_X1    g060(.A(G162gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT79), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(new_n263), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n256), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n254), .A2(KEYINPUT81), .ZN(new_n268));
  OR3_X1    g067(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n254), .A2(KEYINPUT81), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT3), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275));
  INV_X1    g074(.A(new_n266), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(new_n264), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n275), .B(new_n272), .C1(new_n277), .C2(new_n256), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  INV_X1    g078(.A(G113gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(G120gat), .ZN(new_n281));
  INV_X1    g080(.A(G120gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n281), .B(new_n283), .C1(G113gat), .C2(new_n282), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n284), .A2(new_n289), .A3(new_n285), .A4(new_n286), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n280), .A2(G120gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n282), .A2(G113gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n288), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n274), .A2(new_n278), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n267), .A2(new_n273), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT4), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n272), .B1(new_n277), .B2(new_n256), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n299), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n300), .A2(new_n303), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n301), .B2(new_n302), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(new_n299), .A3(KEYINPUT82), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n305), .A2(new_n299), .B1(new_n304), .B2(new_n308), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n307), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n303), .A3(new_n315), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n310), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G57gat), .B(G85gat), .Z(new_n321));
  XNOR2_X1  g120(.A(G1gat), .B(G29gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(KEYINPUT84), .A3(new_n326), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n325), .B(new_n310), .C1(new_n317), .C2(new_n319), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n320), .A2(new_n334), .A3(KEYINPUT6), .A4(new_n326), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT85), .B1(new_n327), .B2(new_n330), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT24), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(G183gat), .A3(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G183gat), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT67), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n204), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(KEYINPUT23), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n204), .A2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n360), .A3(KEYINPUT25), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n339), .B1(new_n351), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n363));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(KEYINPUT23), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n363), .A2(new_n368), .A3(KEYINPUT68), .A4(new_n356), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n344), .B2(new_n347), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n359), .A2(G176gat), .ZN(new_n371));
  OR2_X1    g170(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT65), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n371), .A2(new_n372), .A3(new_n376), .A4(new_n373), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n362), .A2(new_n369), .B1(new_n367), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT27), .B(G183gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n346), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n381), .A2(KEYINPUT28), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n381), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n357), .B1(new_n358), .B2(KEYINPUT26), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n354), .A2(new_n355), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(KEYINPUT26), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n338), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n378), .A2(new_n367), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n356), .A2(new_n360), .A3(KEYINPUT25), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT68), .B1(new_n391), .B2(new_n363), .ZN(new_n392));
  AND4_X1   g191(.A1(KEYINPUT68), .A2(new_n363), .A3(new_n356), .A4(new_n368), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT75), .A3(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n389), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n387), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(KEYINPUT73), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(KEYINPUT73), .B2(new_n404), .ZN(new_n406));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(G64gat), .ZN(new_n412));
  INV_X1    g211(.A(G92gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n379), .A2(new_n338), .A3(new_n388), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT75), .B1(new_n394), .B2(new_n387), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT76), .A3(new_n396), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT76), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n389), .B2(new_n395), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n397), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n399), .A2(new_n397), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n408), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n415), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  AOI211_X1 g227(.A(KEYINPUT77), .B(new_n426), .C1(new_n420), .C2(new_n423), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n410), .B(new_n414), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n414), .A2(KEYINPUT30), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n410), .B(new_n434), .C1(new_n428), .C2(new_n429), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n410), .B1(new_n428), .B2(new_n429), .ZN(new_n436));
  INV_X1    g235(.A(new_n414), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n337), .A2(new_n433), .A3(new_n435), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G22gat), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n408), .B1(new_n278), .B2(new_n400), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT3), .B1(new_n408), .B2(new_n416), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n302), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n408), .A2(new_n400), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n302), .B1(new_n446), .B2(new_n275), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n442), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n440), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n448), .A3(new_n440), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(G50gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n449), .B2(KEYINPUT87), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n452), .B(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n301), .B1(new_n379), .B2(new_n388), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n394), .A2(new_n299), .A3(new_n387), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G43gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n462), .A2(new_n463), .A3(G227gat), .A4(G233gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT72), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT32), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n472), .B2(KEYINPUT32), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n473), .B2(new_n471), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n468), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n468), .A3(new_n480), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n467), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n478), .A2(new_n468), .A3(new_n480), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n485), .A2(new_n481), .A3(new_n466), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n461), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n467), .A3(new_n483), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n466), .B1(new_n485), .B2(new_n481), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT36), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n460), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n409), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n428), .B2(new_n429), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT76), .B1(new_n419), .B2(new_n396), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n422), .A2(new_n421), .A3(new_n397), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n427), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT77), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n424), .A2(new_n415), .A3(new_n427), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n409), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n437), .B(new_n496), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT38), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n327), .A2(new_n330), .A3(new_n332), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n430), .A2(new_n335), .A3(new_n336), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n408), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n424), .A2(new_n509), .A3(new_n425), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n402), .A2(new_n509), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(new_n503), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT38), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n437), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n414), .B1(new_n517), .B2(new_n495), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(KEYINPUT90), .A3(new_n513), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n505), .A2(new_n508), .A3(new_n516), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n458), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n300), .A2(new_n303), .A3(new_n306), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n308), .ZN(new_n523));
  INV_X1    g322(.A(new_n314), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n307), .B1(new_n305), .B2(new_n299), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(KEYINPUT39), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n526), .B(new_n325), .C1(KEYINPUT39), .C2(new_n523), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n327), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n435), .B1(new_n502), .B2(new_n414), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n431), .B1(new_n502), .B2(new_n414), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT88), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n433), .A2(new_n438), .A3(new_n535), .A4(new_n435), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n531), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n493), .B1(new_n521), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n533), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n484), .A2(new_n486), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(new_n337), .A3(new_n458), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n336), .A2(new_n335), .A3(new_n506), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n458), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n484), .B2(new_n486), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT91), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n536), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n253), .B1(new_n538), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G64gat), .Z(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT97), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT96), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n563), .B1(new_n562), .B2(KEYINPUT96), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n554), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n238), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n572), .A2(new_n574), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n576), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n570), .A2(new_n571), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT8), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n597), .C1(G85gat), .C2(G92gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n237), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n600), .A2(new_n232), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT101), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n607), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n610), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT103), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n584), .A2(new_n592), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G230gat), .ZN(new_n622));
  INV_X1    g421(.A(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n565), .A2(new_n566), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n601), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n600), .B1(new_n567), .B2(new_n569), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n570), .A2(new_n601), .A3(new_n629), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n624), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n628), .A2(new_n622), .A3(new_n623), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G176gat), .ZN(new_n636));
  INV_X1    g435(.A(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n633), .B2(new_n634), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n621), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n553), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n337), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n551), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n551), .A4(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n553), .A2(new_n643), .ZN(new_n653));
  INV_X1    g452(.A(new_n551), .ZN(new_n654));
  OAI21_X1  g453(.A(G8gat), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT104), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n651), .A2(new_n655), .A3(new_n658), .A4(new_n652), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n547), .A2(new_n548), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n653), .A2(G15gat), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n491), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(G15gat), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n458), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n593), .A2(new_n620), .ZN(new_n672));
  INV_X1    g471(.A(new_n619), .ZN(new_n673));
  INV_X1    g472(.A(new_n642), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n553), .A2(new_n222), .A3(new_n645), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(new_n531), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n551), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT90), .B1(new_n518), .B2(new_n513), .ZN(new_n681));
  AND4_X1   g480(.A1(KEYINPUT90), .A2(new_n496), .A3(new_n437), .A4(new_n513), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n507), .B1(new_n504), .B2(KEYINPUT38), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n459), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n492), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n654), .A2(new_n549), .B1(new_n541), .B2(KEYINPUT35), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT107), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n538), .A2(new_n552), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n619), .A2(KEYINPUT44), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n673), .B1(new_n686), .B2(new_n687), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n672), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(new_n253), .A3(new_n642), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n696), .A2(new_n337), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n678), .B1(new_n702), .B2(new_n222), .ZN(G1328gat));
  NAND4_X1  g502(.A1(new_n553), .A2(new_n223), .A3(new_n551), .A4(new_n676), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT46), .Z(new_n705));
  NOR3_X1   g504(.A1(new_n696), .A2(new_n654), .A3(new_n701), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n223), .ZN(G1329gat));
  XNOR2_X1  g506(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n695), .A2(new_n664), .A3(new_n700), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n675), .A2(G43gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n553), .A2(new_n661), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n708), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n708), .ZN(new_n714));
  INV_X1    g513(.A(new_n712), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n714), .B(new_n715), .C1(new_n709), .C2(G43gat), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(G1330gat));
  NAND3_X1  g516(.A1(new_n695), .A2(new_n459), .A3(new_n700), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G50gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n675), .A2(G50gat), .A3(new_n458), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n553), .A2(KEYINPUT110), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n553), .A2(new_n720), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n723), .B(KEYINPUT109), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n718), .B2(G50gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g528(.A1(new_n688), .A2(new_n690), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n253), .A2(new_n642), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n621), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n645), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n551), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n733), .B2(new_n491), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n662), .A2(G71gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(new_n732), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n741), .A2(KEYINPUT50), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n734), .A2(new_n459), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g549(.A1(new_n337), .A2(G85gat), .A3(new_n674), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n538), .A2(new_n552), .ZN(new_n752));
  INV_X1    g551(.A(new_n672), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n252), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n673), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n673), .A4(new_n754), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(KEYINPUT112), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT112), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n751), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n753), .A2(new_n731), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n695), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT111), .B1(new_n763), .B2(new_n337), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G85gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n763), .A2(KEYINPUT111), .A3(new_n337), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(G1336gat));
  NAND3_X1  g566(.A1(new_n695), .A2(new_n551), .A3(new_n762), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n758), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n551), .A2(new_n413), .A3(new_n642), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT113), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n776));
  NAND2_X1  g575(.A1(new_n755), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n758), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n768), .A2(G92gat), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  NOR3_X1   g580(.A1(new_n662), .A2(G99gat), .A3(new_n674), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n784), .B(new_n785), .C1(new_n759), .C2(new_n760), .ZN(new_n786));
  OAI21_X1  g585(.A(G99gat), .B1(new_n763), .B2(new_n491), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n695), .A2(new_n459), .A3(new_n762), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n458), .A2(new_n674), .A3(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT53), .B1(new_n770), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n789), .A2(G106gat), .B1(new_n778), .B2(new_n791), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n621), .A2(new_n252), .A3(new_n642), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n638), .B1(new_n633), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n630), .A2(new_n632), .A3(new_n624), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT10), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n803), .A2(new_n631), .B1(new_n622), .B2(new_n623), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT54), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n640), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT117), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n801), .A2(new_n805), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n640), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n808), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n248), .A2(new_n234), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n233), .A2(new_n235), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n206), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n251), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n619), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n808), .A2(new_n252), .A3(new_n811), .A4(new_n813), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n674), .A2(new_n818), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n673), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n698), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n459), .B1(new_n799), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n662), .A2(new_n551), .A3(new_n337), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n280), .A3(new_n253), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n799), .A2(new_n826), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n645), .A3(new_n654), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n832), .A2(new_n459), .A3(new_n486), .A4(new_n484), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n252), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n834), .B2(new_n280), .ZN(G1340gat));
  NOR3_X1   g634(.A1(new_n829), .A2(new_n282), .A3(new_n674), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n642), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n282), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n833), .B2(new_n753), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n827), .A2(G127gat), .A3(new_n699), .A4(new_n828), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n833), .A2(new_n844), .A3(new_n673), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n829), .B2(new_n619), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G1343gat));
  INV_X1    g648(.A(G141gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n664), .A2(new_n551), .A3(new_n337), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT119), .B1(new_n809), .B2(new_n810), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n855), .B(KEYINPUT55), .C1(new_n801), .C2(new_n805), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n252), .A2(new_n640), .A3(new_n806), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n824), .B(KEYINPUT120), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n858), .A2(new_n854), .A3(new_n856), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n823), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n862), .A3(new_n619), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n753), .B1(new_n863), .B2(new_n820), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n799), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n458), .B1(new_n799), .B2(new_n826), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n852), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n850), .B1(new_n871), .B2(new_n252), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n832), .A2(new_n458), .A3(new_n664), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n253), .A2(G141gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT58), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n253), .B(new_n852), .C1(new_n868), .C2(new_n870), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n875), .B(new_n878), .C1(new_n879), .C2(new_n850), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n873), .A2(new_n882), .A3(new_n642), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n882), .C1(new_n871), .C2(new_n642), .ZN(new_n884));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n864), .A2(new_n797), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n459), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n831), .A2(new_n853), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n642), .B(new_n851), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n884), .B2(new_n890), .ZN(G1345gat));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n261), .A3(new_n753), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n871), .A2(new_n699), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n261), .ZN(G1346gat));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n262), .A3(new_n673), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n871), .A2(new_n673), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n262), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n654), .A2(new_n645), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n458), .A2(new_n831), .A3(new_n540), .A4(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n899), .A2(new_n372), .A3(new_n373), .A4(new_n252), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n654), .A2(new_n662), .A3(new_n645), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n827), .A2(KEYINPUT123), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT123), .B1(new_n827), .B2(new_n901), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n902), .A2(new_n903), .A3(new_n253), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n904), .B2(new_n204), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n899), .A2(new_n353), .A3(new_n642), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n902), .A2(new_n903), .A3(new_n674), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n353), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n902), .A2(new_n903), .A3(new_n698), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n345), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n899), .A2(new_n380), .A3(new_n753), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT60), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n915), .B(new_n916), .C1(new_n345), .C2(new_n909), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n346), .A3(new_n673), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n902), .A2(new_n903), .A3(new_n619), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n346), .B1(new_n921), .B2(KEYINPUT61), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(KEYINPUT61), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n920), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  NOR3_X1   g725(.A1(new_n654), .A2(new_n664), .A3(new_n645), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n869), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n252), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n887), .A2(new_n888), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n927), .B(KEYINPUT126), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n252), .A2(G197gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n637), .A3(new_n642), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  NOR3_X1   g735(.A1(new_n930), .A2(new_n674), .A3(new_n931), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n637), .ZN(G1353gat));
  INV_X1    g737(.A(G211gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n939), .A3(new_n753), .ZN(new_n940));
  INV_X1    g739(.A(new_n931), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n753), .B(new_n941), .C1(new_n887), .C2(new_n888), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n928), .B2(new_n673), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n673), .A2(G218gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n932), .B2(new_n948), .ZN(G1355gat));
endmodule


