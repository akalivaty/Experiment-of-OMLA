//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039;
  INV_X1    g000(.A(KEYINPUT21), .ZN(new_n202));
  INV_X1    g001(.A(G71gat), .ZN(new_n203));
  INV_X1    g002(.A(G78gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT97), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(G57gat), .A2(G64gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G57gat), .A2(G64gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(KEYINPUT97), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n207), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT9), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n212), .A3(new_n213), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n202), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(G127gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G22gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G15gat), .ZN(new_n226));
  INV_X1    g025(.A(G15gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G22gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT91), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(KEYINPUT92), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(KEYINPUT92), .B2(new_n232), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n226), .A2(new_n228), .A3(new_n235), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n235), .B1(new_n226), .B2(new_n228), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G8gat), .ZN(new_n242));
  INV_X1    g041(.A(G8gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n215), .A2(new_n219), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(KEYINPUT21), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT98), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT98), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n247), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n223), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G155gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G183gat), .B(G211gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n249), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n249), .B2(new_n252), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261));
  INV_X1    g060(.A(G85gat), .ZN(new_n262));
  INV_X1    g061(.A(G92gat), .ZN(new_n263));
  AOI22_X1  g062(.A1(KEYINPUT8), .A2(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G99gat), .B(G106gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n264), .A2(new_n265), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n270), .A2(new_n218), .ZN(new_n271));
  AND2_X1   g070(.A1(G57gat), .A2(G64gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(G57gat), .A2(G64gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n210), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n214), .A2(new_n274), .A3(KEYINPUT9), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n206), .A3(new_n205), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT8), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n263), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(new_n268), .A3(new_n278), .A4(new_n269), .ZN(new_n279));
  INV_X1    g078(.A(new_n265), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT101), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(KEYINPUT101), .A3(new_n280), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n271), .A2(new_n276), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n270), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(new_n215), .B2(new_n219), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n260), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G120gat), .B(G148gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT103), .ZN(new_n291));
  XNOR2_X1  g090(.A(G176gat), .B(G204gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n260), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT10), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n285), .A2(new_n297), .A3(new_n287), .ZN(new_n298));
  INV_X1    g097(.A(new_n286), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n246), .A2(KEYINPUT10), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT102), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n296), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(KEYINPUT102), .A3(new_n300), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n295), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n296), .B1(new_n298), .B2(new_n300), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n307), .A2(new_n288), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT104), .B1(new_n308), .B2(new_n293), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT104), .B(new_n293), .C1(new_n307), .C2(new_n288), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n306), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G29gat), .ZN(new_n314));
  INV_X1    g113(.A(G36gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT14), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT14), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G29gat), .B2(G36gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(G43gat), .A2(G50gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT15), .ZN(new_n322));
  NAND2_X1  g121(.A1(G43gat), .A2(G50gat), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n321), .A2(KEYINPUT90), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT89), .B(G29gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n320), .B(new_n324), .C1(new_n315), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT15), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n325), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n319), .B1(new_n330), .B2(G36gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(KEYINPUT90), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n299), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT99), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(KEYINPUT99), .A3(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n329), .A2(new_n334), .A3(KEYINPUT17), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT17), .B1(new_n329), .B2(new_n334), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n286), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G134gat), .B(G162gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G190gat), .B(G218gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT100), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n346), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n335), .A2(KEYINPUT99), .A3(new_n336), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT99), .B1(new_n335), .B2(new_n336), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n344), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n351), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n341), .B2(new_n344), .ZN(new_n358));
  INV_X1    g157(.A(new_n355), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n259), .A2(new_n313), .A3(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT73), .ZN(new_n365));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G211gat), .B(G218gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT71), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(G197gat), .A2(G204gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT22), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n372), .A2(new_n373), .B1(new_n376), .B2(new_n375), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n380), .A2(new_n370), .A3(new_n369), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(G183gat), .A3(G190gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT24), .ZN(new_n389));
  NOR2_X1   g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n385), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n384), .A2(G169gat), .A3(G176gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G169gat), .ZN(new_n399));
  INV_X1    g198(.A(G176gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT65), .B(new_n396), .C1(new_n401), .C2(new_n384), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n393), .A2(KEYINPUT66), .A3(new_n398), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT66), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n402), .ZN(new_n405));
  OR2_X1    g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT24), .A3(new_n388), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n407), .A2(KEYINPUT25), .A3(new_n385), .A4(new_n387), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n396), .B1(new_n401), .B2(new_n384), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n392), .B1(new_n391), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT64), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT64), .B(new_n392), .C1(new_n391), .C2(new_n410), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n403), .A2(new_n409), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT27), .B(G183gat), .ZN(new_n416));
  INV_X1    g215(.A(G190gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OR3_X1    g217(.A1(new_n418), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n419));
  XOR2_X1   g218(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n401), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n422), .A2(KEYINPUT26), .A3(new_n397), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n422), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n419), .A2(new_n421), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n415), .A2(new_n425), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n383), .B(new_n427), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n415), .A2(new_n425), .A3(new_n426), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n415), .B2(new_n425), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n382), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT72), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n431), .A2(new_n432), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT72), .A3(new_n383), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n368), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n437), .A3(new_n368), .ZN(new_n440));
  AND2_X1   g239(.A1(KEYINPUT74), .A2(KEYINPUT30), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(KEYINPUT74), .A2(KEYINPUT30), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n368), .B(new_n445), .C1(new_n435), .C2(new_n437), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n453));
  INV_X1    g252(.A(G141gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G148gat), .ZN(new_n455));
  INV_X1    g254(.A(G148gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G141gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT76), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G155gat), .B(G162gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(G162gat), .ZN(new_n465));
  INV_X1    g264(.A(G162gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(KEYINPUT77), .ZN(new_n467));
  OAI21_X1  g266(.A(G155gat), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT78), .B1(new_n468), .B2(KEYINPUT2), .ZN(new_n469));
  INV_X1    g268(.A(G155gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(KEYINPUT77), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(G162gat), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT78), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT2), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n463), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n470), .A2(new_n466), .A3(KEYINPUT75), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT75), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(G155gat), .B2(G162gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT2), .B1(new_n455), .B2(new_n457), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n477), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G127gat), .B(G134gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G113gat), .B(G120gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(KEYINPUT1), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT1), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT80), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT77), .B(G162gat), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT78), .B(KEYINPUT2), .C1(new_n501), .C2(new_n470), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n462), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT79), .B1(new_n503), .B2(new_n485), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n491), .A2(new_n494), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n477), .A2(new_n486), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n453), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n487), .A2(new_n504), .A3(KEYINPUT3), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n500), .A2(new_n502), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n485), .B1(new_n513), .B2(new_n463), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT3), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n514), .A2(new_n515), .B1(new_n497), .B2(new_n498), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n510), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n477), .A2(new_n518), .A3(new_n486), .A4(new_n506), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n514), .A2(KEYINPUT81), .A3(new_n518), .A4(new_n506), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n511), .A2(new_n525), .ZN(new_n526));
  AOI211_X1 g325(.A(KEYINPUT5), .B(new_n510), .C1(new_n512), .C2(new_n516), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT82), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n514), .A2(KEYINPUT82), .A3(new_n518), .A4(new_n506), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n523), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT83), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  AND4_X1   g331(.A1(KEYINPUT83), .A2(new_n517), .A3(new_n453), .A4(new_n531), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n452), .B(new_n526), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n453), .A3(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT83), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n527), .A2(KEYINPUT83), .A3(new_n531), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n452), .B1(new_n541), .B2(new_n526), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n544));
  INV_X1    g343(.A(new_n452), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT6), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n448), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n415), .A2(new_n506), .A3(new_n425), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n506), .B1(new_n415), .B2(new_n425), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT33), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(KEYINPUT32), .ZN(new_n556));
  XOR2_X1   g355(.A(G15gat), .B(G43gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT68), .ZN(new_n558));
  XNOR2_X1  g357(.A(G71gat), .B(G99gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n415), .A2(new_n425), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n495), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n415), .A2(new_n506), .A3(new_n425), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n566), .B2(new_n550), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(KEYINPUT33), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT69), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n553), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n568), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n561), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n549), .A3(new_n565), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT34), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n553), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n570), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n574), .A3(new_n561), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n503), .A2(KEYINPUT3), .A3(new_n485), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n382), .B1(new_n582), .B2(KEYINPUT29), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n379), .B2(new_n381), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n515), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n487), .A2(new_n586), .A3(new_n504), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G228gat), .ZN(new_n589));
  INV_X1    g388(.A(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n378), .A2(new_n369), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT29), .B1(new_n378), .B2(new_n369), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT3), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n593), .B1(new_n514), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n583), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n592), .A2(new_n225), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n593), .B1(new_n583), .B2(new_n587), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n514), .A2(new_n515), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n584), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n603), .B2(new_n382), .ZN(new_n604));
  OAI21_X1  g403(.A(G22gat), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT84), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G78gat), .B(G106gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n588), .A2(new_n591), .B1(new_n583), .B2(new_n598), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT84), .B1(new_n611), .B2(new_n225), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n605), .A3(new_n608), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT31), .B(G50gat), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n610), .B2(new_n613), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n576), .B(new_n581), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT35), .B1(new_n548), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n580), .A2(new_n574), .A3(new_n561), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n574), .B1(new_n580), .B2(new_n561), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n581), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n614), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n608), .B1(new_n612), .B2(new_n605), .ZN(new_n626));
  AND4_X1   g425(.A1(new_n606), .A2(new_n600), .A3(new_n605), .A4(new_n608), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n544), .A2(new_n545), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(new_n535), .A3(new_n534), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n632), .A2(new_n546), .B1(new_n442), .B2(new_n447), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n624), .A2(new_n630), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n616), .ZN(new_n636));
  NOR2_X1   g435(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT70), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n576), .B(new_n581), .C1(new_n637), .C2(new_n640), .ZN(new_n641));
  OAI22_X1  g440(.A1(new_n620), .A2(new_n621), .B1(new_n638), .B2(new_n639), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n548), .A2(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n435), .A2(new_n437), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n367), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n435), .A2(KEYINPUT37), .A3(new_n437), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT38), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n430), .A2(new_n433), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT38), .B1(new_n650), .B2(KEYINPUT37), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n438), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n649), .A2(new_n632), .A3(new_n546), .A4(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n440), .A2(new_n441), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n446), .B1(new_n654), .B2(new_n439), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT85), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n512), .A2(new_n516), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n509), .B1(new_n531), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n452), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT39), .B1(new_n508), .B2(new_n510), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n656), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n656), .B(new_n666), .C1(new_n661), .C2(new_n663), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n655), .A2(new_n631), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n668), .A3(new_n630), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n618), .A2(new_n635), .B1(new_n643), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G169gat), .B(G197gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT12), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n237), .A2(new_n240), .A3(new_n243), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n243), .B1(new_n237), .B2(new_n240), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n680), .B(KEYINPUT93), .C1(new_n342), .C2(new_n343), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n329), .A2(new_n334), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT17), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n329), .A2(new_n334), .A3(KEYINPUT17), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n245), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT93), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n680), .B2(new_n682), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n681), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G229gat), .A2(G233gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(KEYINPUT18), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n245), .B(new_n682), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n691), .B(KEYINPUT13), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n689), .B2(new_n691), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n677), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n689), .A2(new_n691), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n697), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n702), .A2(new_n692), .A3(new_n695), .A4(new_n676), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT96), .B1(new_n670), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n635), .A2(new_n618), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n548), .A2(new_n636), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n641), .A2(new_n642), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n669), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT96), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n704), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n363), .B1(new_n706), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n632), .A2(new_n546), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g517(.A(KEYINPUT16), .B(G8gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n714), .A2(new_n655), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n243), .B1(new_n714), .B2(new_n655), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT42), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n714), .A2(new_n655), .A3(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(G1325gat));
  AOI21_X1  g526(.A(G15gat), .B1(new_n714), .B2(new_n624), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n709), .A2(new_n227), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT105), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n714), .B2(new_n730), .ZN(G1326gat));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n636), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  INV_X1    g533(.A(new_n259), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n313), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n362), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n706), .B2(new_n713), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n715), .A2(new_n330), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(KEYINPUT45), .A3(new_n740), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n670), .B2(new_n362), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n653), .A2(new_n668), .A3(new_n630), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n640), .A2(new_n637), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n620), .A2(new_n621), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n640), .B1(new_n576), .B2(new_n581), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n633), .A2(new_n630), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n636), .B1(new_n623), .B2(new_n622), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n715), .A2(new_n448), .A3(new_n634), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n620), .A2(new_n621), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n715), .A2(new_n630), .A3(new_n755), .A4(new_n448), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n753), .A2(new_n754), .B1(new_n756), .B2(KEYINPUT35), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT44), .B(new_n361), .C1(new_n752), .C2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n736), .A2(new_n705), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(new_n716), .A3(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n743), .B(new_n744), .C1(new_n761), .C2(new_n325), .ZN(G1328gat));
  NAND2_X1  g561(.A1(new_n706), .A2(new_n713), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n737), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n655), .A2(new_n315), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT46), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n759), .A2(new_n655), .A3(new_n760), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n766), .B(new_n767), .C1(new_n315), .C2(new_n768), .ZN(G1329gat));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  INV_X1    g569(.A(new_n709), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(G43gat), .ZN(new_n772));
  AND4_X1   g571(.A1(new_n746), .A2(new_n758), .A3(new_n760), .A4(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n739), .A2(new_n624), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n770), .B(new_n774), .C1(new_n775), .C2(G43gat), .ZN(new_n776));
  AOI21_X1  g575(.A(G43gat), .B1(new_n739), .B2(new_n624), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT47), .B1(new_n777), .B2(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1330gat));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n636), .A2(G50gat), .ZN(new_n781));
  AND4_X1   g580(.A1(new_n746), .A2(new_n758), .A3(new_n760), .A4(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n739), .A2(new_n636), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n780), .B(new_n783), .C1(new_n784), .C2(G50gat), .ZN(new_n785));
  AOI21_X1  g584(.A(G50gat), .B1(new_n739), .B2(new_n636), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT48), .B1(new_n786), .B2(new_n782), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1331gat));
  NAND3_X1  g587(.A1(new_n259), .A2(new_n362), .A3(new_n312), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n670), .A2(new_n704), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n716), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n655), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT106), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT107), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(KEYINPUT107), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(G1333gat));
  NAND2_X1  g601(.A1(new_n790), .A2(new_n624), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n203), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n709), .A2(new_n203), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n790), .A2(KEYINPUT108), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT108), .B1(new_n790), .B2(new_n805), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n804), .B(new_n809), .C1(new_n806), .C2(new_n807), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1334gat));
  NAND2_X1  g612(.A1(new_n790), .A2(new_n636), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g614(.A1(new_n259), .A2(new_n704), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n361), .B(new_n816), .C1(new_n752), .C2(new_n757), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n362), .B1(new_n707), .B2(new_n710), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n816), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n716), .A2(new_n262), .A3(new_n312), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT110), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n259), .A2(new_n704), .A3(new_n313), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n746), .A2(new_n716), .A3(new_n758), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G85gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT111), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n825), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1336gat));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n655), .A2(new_n263), .A3(new_n312), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT112), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n822), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n746), .A2(new_n655), .A3(new_n758), .A4(new_n826), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G92gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AND4_X1   g642(.A1(KEYINPUT51), .A2(new_n711), .A3(new_n361), .A4(new_n816), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT51), .B1(new_n820), .B2(new_n816), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n839), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n837), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n842), .A2(new_n846), .A3(new_n847), .A4(new_n836), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n843), .A2(new_n848), .ZN(G1337gat));
  NAND3_X1  g648(.A1(new_n759), .A2(new_n771), .A3(new_n826), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G99gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n313), .A2(G99gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n822), .A2(new_n624), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1338gat));
  NOR3_X1   g653(.A1(new_n630), .A2(G106gat), .A3(new_n313), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n822), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n746), .A2(new_n636), .A3(new_n758), .A4(new_n826), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G106gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1339gat));
  INV_X1    g662(.A(new_n753), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n301), .A2(new_n302), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n304), .A3(new_n260), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n298), .A2(new_n300), .A3(new_n296), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT54), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n871), .B(new_n294), .C1(new_n307), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n305), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n868), .B1(new_n303), .B2(new_n304), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n307), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n293), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n871), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n700), .B2(new_n703), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n693), .A2(new_n694), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n689), .B2(new_n691), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n675), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n703), .A2(new_n312), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n362), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n703), .A2(new_n883), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT114), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n874), .A2(new_n878), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n703), .A2(new_n889), .A3(new_n883), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n361), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n259), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n363), .A2(new_n704), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT115), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n704), .A2(new_n888), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n703), .A2(new_n312), .A3(new_n883), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n361), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n703), .A2(new_n889), .A3(new_n883), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n889), .B1(new_n703), .B2(new_n883), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n361), .A2(new_n878), .A3(new_n874), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n735), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n363), .A2(new_n704), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n864), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n715), .A2(new_n655), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G113gat), .B1(new_n908), .B2(new_n705), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n715), .B1(new_n894), .B2(new_n905), .ZN(new_n910));
  INV_X1    g709(.A(new_n617), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n448), .A3(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n705), .A2(G113gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1340gat));
  INV_X1    g715(.A(G120gat), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n908), .A2(new_n917), .A3(new_n313), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n912), .A2(new_n313), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n917), .ZN(G1341gat));
  OAI21_X1  g719(.A(G127gat), .B1(new_n908), .B2(new_n735), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n735), .A2(G127gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n912), .B2(new_n922), .ZN(G1342gat));
  NAND2_X1  g722(.A1(new_n448), .A2(new_n361), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT117), .Z(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(G134gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n928));
  OAI21_X1  g727(.A(G134gat), .B1(new_n908), .B2(new_n362), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(G1343gat));
  NAND2_X1  g730(.A1(new_n894), .A2(new_n905), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n636), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n709), .A2(new_n907), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n636), .B1(new_n892), .B2(new_n893), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(KEYINPUT57), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G141gat), .B1(new_n938), .B2(new_n705), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n709), .A2(new_n636), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n910), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n932), .A2(new_n716), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT118), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n705), .A2(G141gat), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n942), .A2(new_n944), .A3(new_n448), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT58), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT58), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n939), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1344gat));
  NAND2_X1  g750(.A1(new_n942), .A2(new_n944), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n953), .A2(new_n456), .A3(new_n448), .A4(new_n312), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n934), .A2(new_n937), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT59), .B(new_n456), .C1(new_n955), .C2(new_n312), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT59), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n935), .A2(new_n313), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n936), .A2(new_n933), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n636), .A2(KEYINPUT57), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n960), .B1(new_n894), .B2(new_n905), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g762(.A(KEYINPUT119), .B(new_n960), .C1(new_n894), .C2(new_n905), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n957), .B1(new_n965), .B2(G148gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n954), .B1(new_n956), .B2(new_n966), .ZN(G1345gat));
  NAND3_X1  g766(.A1(new_n953), .A2(new_n448), .A3(new_n259), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n259), .A2(G155gat), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT120), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n968), .A2(new_n470), .B1(new_n955), .B2(new_n970), .ZN(G1346gat));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n972));
  INV_X1    g771(.A(new_n925), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n501), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n952), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n501), .B1(new_n955), .B2(new_n361), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n938), .A2(new_n362), .ZN(new_n978));
  OAI221_X1 g777(.A(KEYINPUT121), .B1(new_n952), .B2(new_n974), .C1(new_n978), .C2(new_n501), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1347gat));
  NOR2_X1   g779(.A1(new_n716), .A2(new_n448), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n932), .A2(new_n753), .A3(new_n981), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n982), .A2(new_n399), .A3(new_n705), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n716), .B1(new_n894), .B2(new_n905), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n617), .A2(new_n448), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(new_n704), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n983), .B1(new_n988), .B2(new_n399), .ZN(G1348gat));
  NOR3_X1   g788(.A1(new_n982), .A2(new_n400), .A3(new_n313), .ZN(new_n990));
  AOI21_X1  g789(.A(G176gat), .B1(new_n987), .B2(new_n312), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n991), .A2(KEYINPUT122), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(KEYINPUT122), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1349gat));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n982), .B2(new_n735), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n906), .A2(KEYINPUT123), .A3(new_n259), .A4(new_n981), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n996), .A2(G183gat), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n987), .A2(new_n416), .A3(new_n259), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(KEYINPUT60), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT60), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n998), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1350gat));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n417), .A3(new_n361), .ZN(new_n1005));
  OAI21_X1  g804(.A(G190gat), .B1(new_n982), .B2(new_n362), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1351gat));
  NOR2_X1   g808(.A1(new_n940), .A2(new_n448), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n932), .A2(new_n715), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n984), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n705), .A2(G197gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g815(.A(new_n1016), .B(KEYINPUT125), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n981), .A2(new_n709), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1018), .B1(new_n963), .B2(new_n964), .ZN(new_n1019));
  OAI21_X1  g818(.A(G197gat), .B1(new_n1019), .B2(new_n705), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1017), .A2(new_n1020), .ZN(G1352gat));
  OAI21_X1  g820(.A(G204gat), .B1(new_n1019), .B2(new_n313), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g824(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n312), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1025), .B1(new_n1011), .B2(new_n1027), .ZN(new_n1028));
  OR3_X1    g827(.A1(new_n1011), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n1022), .A2(new_n1028), .A3(new_n1029), .ZN(G1353gat));
  NOR2_X1   g829(.A1(new_n735), .A2(G211gat), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1012), .A2(new_n1014), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g831(.A(new_n259), .B(new_n1018), .C1(new_n963), .C2(new_n964), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1033), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1034));
  AOI21_X1  g833(.A(KEYINPUT63), .B1(new_n1033), .B2(G211gat), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(G1354gat));
  OAI21_X1  g835(.A(G218gat), .B1(new_n1019), .B2(new_n362), .ZN(new_n1037));
  NOR2_X1   g836(.A1(new_n362), .A2(G218gat), .ZN(new_n1038));
  NAND3_X1  g837(.A1(new_n1012), .A2(new_n1014), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1037), .A2(new_n1039), .ZN(G1355gat));
endmodule


