//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g0025(.A1(G87), .A2(G250), .ZN(new_n226));
  NOR4_X1   g0026(.A1(new_n219), .A2(new_n222), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT65), .B(G77), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G244), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n209), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n208), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n213), .B(new_n232), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G150), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(KEYINPUT8), .A3(new_n258), .ZN(new_n259));
  OR3_X1    g0059(.A1(new_n223), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n208), .A2(G33), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT69), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n254), .B1(new_n208), .B2(new_n201), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n233), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n207), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT70), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n208), .A2(G1), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(G13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(new_n233), .A3(new_n266), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n271), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n265), .A2(new_n267), .B1(new_n276), .B2(G50), .ZN(new_n277));
  INV_X1    g0077(.A(new_n274), .ZN(new_n278));
  INV_X1    g0078(.A(G50), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT73), .A3(KEYINPUT9), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n277), .A2(new_n280), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT66), .B(G1698), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n290), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n229), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n295), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n294), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(G200), .B2(new_n300), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n286), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT71), .B(G179), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n300), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n281), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n289), .A2(G238), .A3(new_n295), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT74), .B1(new_n315), .B2(new_n297), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n297), .A3(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n298), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n224), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n292), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n289), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n319), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n315), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n316), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n289), .B1(new_n326), .B2(new_n327), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT13), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n253), .A2(G50), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n217), .A2(G20), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n264), .C2(new_n202), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n267), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n276), .A2(G68), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n270), .A2(new_n273), .A3(new_n217), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT12), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(new_n267), .A3(new_n343), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n345), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n332), .A2(new_n336), .A3(G190), .ZN(new_n352));
  AND4_X1   g0152(.A1(KEYINPUT76), .A2(new_n338), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n337), .B2(G200), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT76), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT77), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n337), .A2(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT14), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n337), .A2(new_n359), .A3(G169), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n358), .B(new_n360), .C1(new_n361), .C2(new_n337), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n350), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n338), .A2(new_n351), .A3(new_n352), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT76), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT77), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n352), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n356), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n297), .B1(new_n299), .B2(new_n224), .ZN(new_n371));
  AND2_X1   g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n375));
  OAI21_X1  g0175(.A(G223), .B1(new_n375), .B2(new_n320), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G226), .A2(G1698), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n329), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT81), .B(new_n329), .C1(new_n378), .C2(new_n380), .ZN(new_n384));
  AOI211_X1 g0184(.A(G190), .B(new_n371), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n371), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT82), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n292), .A2(new_n392), .A3(G20), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n374), .B2(new_n208), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n255), .A2(G58), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n258), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n398), .B2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT78), .B1(new_n399), .B2(new_n208), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT67), .B(G58), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n217), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n401), .B(G20), .C1(new_n403), .C2(new_n396), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n253), .A2(G159), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n395), .A2(new_n400), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n392), .B1(new_n292), .B2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(G68), .B1(G159), .B2(new_n253), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n400), .A4(new_n404), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n413), .A3(new_n267), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n261), .B2(new_n268), .ZN(new_n416));
  AOI211_X1 g0216(.A(KEYINPUT79), .B(new_n271), .C1(new_n259), .C2(new_n260), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n416), .A2(new_n417), .A3(new_n275), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT80), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n261), .A2(new_n274), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n261), .A2(new_n268), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n267), .B1(new_n270), .B2(new_n273), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n261), .A2(new_n415), .A3(new_n268), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n420), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT80), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n290), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n379), .B1(new_n430), .B2(new_n374), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT81), .B1(new_n431), .B2(new_n329), .ZN(new_n432));
  INV_X1    g0232(.A(new_n384), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n301), .B(new_n386), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT82), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n389), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n391), .A2(new_n414), .A3(new_n429), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(KEYINPUT83), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(KEYINPUT83), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n408), .A2(new_n413), .A3(new_n267), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n426), .A2(KEYINPUT80), .A3(new_n427), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(new_n440), .A3(new_n391), .A4(new_n436), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n309), .B1(new_n383), .B2(new_n384), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n386), .B1(new_n311), .B2(new_n387), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n444), .B2(new_n447), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n414), .A2(new_n445), .A3(new_n446), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT18), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n375), .A2(new_n320), .ZN(new_n459));
  OAI221_X1 g0259(.A(new_n292), .B1(new_n218), .B2(new_n324), .C1(new_n459), .C2(new_n224), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n329), .C1(G107), .C2(new_n292), .ZN(new_n461));
  INV_X1    g0261(.A(new_n299), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G244), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n297), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n309), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT15), .B(G87), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n263), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT72), .ZN(new_n468));
  INV_X1    g0268(.A(new_n253), .ZN(new_n469));
  XOR2_X1   g0269(.A(KEYINPUT8), .B(G58), .Z(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI221_X1 g0271(.A(new_n468), .B1(new_n208), .B2(new_n228), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n267), .B1(G77), .B2(new_n276), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n278), .A2(new_n228), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n464), .A2(new_n311), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n450), .A2(new_n458), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n474), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n464), .A2(new_n301), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n464), .A2(G200), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NOR4_X1   g0282(.A1(new_n314), .A2(new_n370), .A3(new_n478), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n411), .A2(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n469), .A2(new_n202), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n220), .A2(new_n487), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n204), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G20), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n484), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n267), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n278), .A2(new_n220), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT84), .B1(new_n287), .B2(G1), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n287), .A2(KEYINPUT84), .A3(G1), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n424), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G97), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G1), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n288), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G41), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .A4(G274), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n289), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(new_n221), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  OAI21_X1  g0311(.A(G244), .B1(new_n375), .B2(new_n320), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n374), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n292), .A2(new_n290), .A3(KEYINPUT4), .A4(G244), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(new_n329), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n518), .A2(G169), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n329), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n521));
  INV_X1    g0321(.A(new_n309), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n507), .C1(new_n509), .C2(new_n221), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n501), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n493), .A2(new_n267), .B1(new_n220), .B2(new_n278), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n518), .A2(G190), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n500), .A4(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n292), .A2(new_n290), .A3(G250), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G294), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n509), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n536), .A2(new_n329), .B1(new_n537), .B2(G264), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n507), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT89), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(KEYINPUT89), .A3(new_n507), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n301), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(new_n388), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n208), .B(G87), .C1(new_n372), .C2(new_n373), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n292), .A2(new_n548), .A3(new_n208), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n208), .A2(G107), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT23), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n550), .A2(KEYINPUT24), .A3(new_n551), .A4(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n267), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n270), .A2(new_n273), .A3(new_n487), .ZN(new_n559));
  NOR2_X1   g0359(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n562));
  INV_X1    g0362(.A(new_n560), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n270), .A2(new_n273), .A3(new_n487), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT88), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n424), .A2(G107), .A3(new_n496), .A4(new_n497), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n558), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n545), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n311), .B1(new_n541), .B2(new_n542), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n539), .A2(new_n361), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n532), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n266), .A2(new_n233), .B1(G20), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n515), .B(new_n208), .C1(G33), .C2(new_n220), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n580), .A2(KEYINPUT20), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT20), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n582), .A2(new_n583), .B1(G116), .B2(new_n274), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n499), .B2(G116), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n537), .A2(G270), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n292), .B(new_n587), .C1(new_n459), .C2(new_n221), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n374), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n329), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(new_n591), .A3(new_n507), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n578), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n278), .A2(new_n579), .ZN(new_n595));
  OAI221_X1 g0395(.A(new_n595), .B1(new_n583), .B2(new_n582), .C1(new_n498), .C2(new_n579), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT21), .A3(G169), .A4(new_n592), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n592), .A2(new_n361), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n596), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT86), .ZN(new_n602));
  OAI21_X1  g0402(.A(G238), .B1(new_n375), .B2(new_n320), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G244), .A2(G1698), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n374), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n287), .A2(new_n579), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n329), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n503), .A2(G274), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n289), .B(G250), .C1(G1), .C2(new_n502), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G200), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n424), .A2(G87), .A3(new_n496), .A4(new_n497), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n292), .A2(new_n208), .A3(G68), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n208), .B1(new_n327), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(G87), .B2(new_n205), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n263), .B2(new_n220), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n267), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n278), .A2(new_n466), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n612), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n607), .A2(G190), .A3(new_n608), .A4(new_n609), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n611), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n610), .A2(new_n311), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n607), .A2(new_n522), .A3(new_n608), .A4(new_n609), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n619), .B(new_n620), .C1(new_n498), .C2(new_n466), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n602), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n623), .A2(new_n627), .A3(new_n602), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n592), .A2(G200), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n585), .B(new_n631), .C1(new_n301), .C2(new_n592), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n601), .A2(new_n629), .A3(new_n630), .A4(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n577), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n483), .A2(new_n634), .ZN(G372));
  INV_X1    g0435(.A(KEYINPUT91), .ZN(new_n636));
  INV_X1    g0436(.A(new_n542), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT89), .B1(new_n538), .B2(new_n507), .ZN(new_n638));
  OAI21_X1  g0438(.A(G169), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n575), .ZN(new_n640));
  INV_X1    g0440(.A(new_n570), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n568), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n639), .A2(new_n640), .B1(new_n642), .B2(new_n558), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n636), .B1(new_n643), .B2(new_n600), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n571), .B1(new_n543), .B2(new_n544), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n526), .A2(new_n531), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n601), .A2(new_n576), .A3(KEYINPUT91), .ZN(new_n648));
  INV_X1    g0448(.A(new_n627), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n621), .A2(new_n622), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n610), .B2(G200), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n610), .A2(new_n651), .A3(G200), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n644), .A2(new_n647), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n526), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT26), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n629), .A2(new_n657), .A3(new_n630), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n656), .A2(new_n659), .A3(new_n627), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n483), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT92), .ZN(new_n664));
  INV_X1    g0464(.A(new_n313), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n477), .B1(new_n366), .B2(new_n368), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n350), .B2(new_n362), .ZN(new_n667));
  INV_X1    g0467(.A(new_n450), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n458), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n669), .B2(new_n308), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(G369));
  NOR2_X1   g0471(.A1(new_n269), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n207), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n596), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n600), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT94), .Z(new_n682));
  NAND4_X1  g0482(.A1(new_n632), .A2(new_n594), .A3(new_n597), .A4(new_n599), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT95), .ZN(new_n687));
  INV_X1    g0487(.A(new_n678), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n572), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n571), .A2(KEYINPUT95), .A3(new_n678), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n573), .A3(new_n576), .A4(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n576), .B2(new_n688), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n576), .A2(new_n678), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n600), .A2(new_n688), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n211), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n235), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n662), .A2(new_n688), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT98), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n532), .A2(new_n573), .A3(new_n655), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n643), .A2(new_n600), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n601), .A2(new_n576), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n647), .A2(new_n714), .A3(KEYINPUT98), .A4(new_n655), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n649), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n712), .A2(new_n713), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n688), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n708), .B1(new_n707), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT96), .B(KEYINPUT30), .Z(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n598), .A2(new_n518), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n536), .A2(new_n329), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n537), .A2(G264), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(new_n610), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n721), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(new_n610), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n598), .A4(new_n518), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n309), .B1(new_n538), .B2(new_n507), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n527), .A3(new_n610), .A4(new_n592), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n678), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n630), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(new_n683), .A3(new_n628), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n647), .A3(new_n576), .A4(new_n688), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n737), .B2(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n727), .A2(new_n731), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(KEYINPUT97), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n729), .B1(new_n739), .B2(KEYINPUT97), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT31), .B(new_n678), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(G330), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n719), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n705), .B1(new_n745), .B2(G1), .ZN(G364));
  OR2_X1    g0546(.A1(new_n684), .A2(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n672), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n701), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n685), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n208), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n292), .B1(new_n754), .B2(G329), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n309), .A2(new_n751), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n388), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(KEYINPUT33), .B(G317), .Z(new_n759));
  OAI21_X1  g0559(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n756), .A2(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n301), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n208), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n762), .A2(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n208), .A2(new_n301), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n309), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n388), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G326), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT100), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n388), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n751), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n760), .B(new_n772), .C1(G283), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n773), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n589), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n769), .A2(G200), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G322), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT101), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n762), .A2(new_n228), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n754), .A2(G159), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  INV_X1    g0584(.A(new_n779), .ZN(new_n785));
  INV_X1    g0585(.A(new_n770), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n292), .B1(new_n785), .B2(new_n402), .C1(new_n279), .C2(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n784), .B(new_n787), .C1(G68), .C2(new_n757), .ZN(new_n788));
  INV_X1    g0588(.A(new_n777), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G87), .A2(new_n789), .B1(new_n775), .B2(G107), .ZN(new_n790));
  INV_X1    g0590(.A(new_n765), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G97), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n781), .B1(new_n782), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n233), .B1(G20), .B2(new_n311), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n795), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n211), .A2(new_n292), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G355), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n699), .A2(new_n292), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n236), .A2(new_n502), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(new_n251), .C2(new_n502), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(G116), .C2(new_n211), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n794), .A2(new_n795), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n684), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n750), .B1(new_n809), .B2(new_n749), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n477), .A2(new_n678), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n688), .B1(new_n473), .B2(new_n474), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n482), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n813), .B2(new_n477), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n706), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(new_n744), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n749), .ZN(new_n817));
  INV_X1    g0617(.A(new_n814), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n796), .ZN(new_n819));
  INV_X1    g0619(.A(new_n749), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n792), .B(new_n374), .C1(new_n763), .C2(new_n753), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G116), .A2(new_n761), .B1(new_n757), .B2(G283), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n823), .B2(KEYINPUT103), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n789), .A2(G107), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT103), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n822), .A2(new_n826), .B1(G294), .B2(new_n779), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n770), .A2(G303), .B1(G87), .B2(new_n775), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G143), .A2(new_n779), .B1(new_n761), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n786), .C1(new_n832), .C2(new_n758), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT34), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n753), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n774), .A2(new_n217), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G50), .C2(new_n789), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n292), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n765), .A2(new_n402), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n829), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n795), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n795), .A2(new_n796), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT102), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n202), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n819), .A2(new_n820), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n817), .A2(new_n846), .ZN(G384));
  NAND3_X1  g0647(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT110), .Z(new_n849));
  INV_X1    g0649(.A(KEYINPUT31), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n634), .B2(new_n688), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n851), .B2(new_n734), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n483), .A2(G330), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n434), .A2(new_n435), .A3(new_n389), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n435), .B1(new_n434), .B2(new_n389), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n856), .A2(new_n448), .B1(new_n441), .B2(new_n440), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n456), .A2(new_n854), .A3(new_n855), .A4(new_n439), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n458), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n676), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n414), .A2(new_n427), .A3(new_n426), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n451), .A2(new_n386), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n387), .A2(new_n311), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n414), .B2(new_n429), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT37), .B1(new_n866), .B2(KEYINPUT106), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n456), .A2(new_n860), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT106), .B1(new_n456), .B2(new_n452), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n867), .A2(new_n437), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n861), .B1(new_n452), .B2(new_n860), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n437), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n437), .A2(new_n868), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n869), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n437), .A2(new_n453), .A3(new_n868), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(new_n867), .B1(KEYINPUT37), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT108), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n857), .B2(new_n858), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n443), .A2(KEYINPUT108), .A3(new_n449), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n458), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n868), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n876), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n848), .B(KEYINPUT110), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n733), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n351), .A2(new_n688), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n366), .B2(new_n368), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n370), .A2(new_n893), .B1(new_n363), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n892), .A2(new_n895), .A3(new_n818), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n862), .A2(new_n875), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT40), .B1(new_n900), .B2(new_n876), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n897), .A2(KEYINPUT40), .B1(new_n901), .B2(new_n896), .ZN(new_n902));
  INV_X1    g0702(.A(G330), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n853), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n883), .A2(new_n458), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT108), .B1(new_n443), .B2(new_n449), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n885), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n880), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n676), .B1(new_n450), .B2(new_n458), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n910), .A2(new_n861), .B1(new_n874), .B2(new_n871), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n909), .A2(new_n887), .B1(KEYINPUT38), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n370), .A2(new_n893), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n894), .A2(new_n363), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n852), .A2(new_n814), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT40), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n901), .A2(new_n896), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n483), .A3(new_n852), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n904), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n662), .A2(new_n814), .A3(new_n688), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n811), .B(KEYINPUT105), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n895), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n862), .B2(new_n875), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n925), .A2(new_n928), .B1(new_n458), .B2(new_n860), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n363), .A2(new_n678), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT39), .B1(new_n926), .B2(new_n927), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n933), .B(new_n876), .C1(new_n886), .C2(new_n888), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n921), .B(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n708), .B(new_n483), .C1(new_n707), .C2(new_n718), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n670), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT109), .Z(new_n941));
  XNOR2_X1  g0741(.A(new_n938), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n207), .B2(new_n672), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n403), .A2(new_n235), .A3(new_n228), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n217), .A2(G50), .ZN(new_n945));
  OAI211_X1 g0745(.A(G1), .B(new_n269), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n579), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n947), .B(new_n234), .C1(KEYINPUT35), .C2(new_n491), .ZN(new_n948));
  XOR2_X1   g0748(.A(KEYINPUT104), .B(KEYINPUT36), .Z(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n946), .A3(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n697), .A2(new_n695), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n646), .B1(new_n501), .B2(new_n678), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n695), .A2(KEYINPUT42), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT42), .B1(new_n697), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n526), .C2(new_n678), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT43), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n655), .B1(new_n621), .B2(new_n688), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n627), .A2(new_n621), .A3(new_n688), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n958), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n959), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n693), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n657), .A2(new_n678), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n956), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n966), .B(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n700), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n969), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n952), .B(new_n973), .C1(KEYINPUT111), .C2(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g0774(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n697), .A2(new_n969), .A3(new_n695), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT45), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n967), .ZN(new_n980));
  INV_X1    g0780(.A(new_n696), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n697), .B1(new_n692), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n685), .B2(KEYINPUT112), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n685), .A2(KEYINPUT112), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n983), .B(new_n984), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n745), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n987), .B2(new_n745), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n748), .A2(G1), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n971), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n766), .A2(new_n758), .B1(new_n786), .B2(new_n763), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n292), .B(new_n991), .C1(G303), .C2(new_n779), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n777), .A2(new_n579), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n993), .A2(KEYINPUT46), .B1(new_n487), .B2(new_n765), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n220), .B2(new_n774), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G317), .C2(new_n754), .ZN(new_n997));
  INV_X1    g0797(.A(G283), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n992), .B(new_n997), .C1(new_n998), .C2(new_n762), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n770), .A2(G143), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n762), .B2(new_n279), .C1(new_n832), .C2(new_n785), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n791), .A2(G68), .ZN(new_n1002));
  INV_X1    g0802(.A(G159), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n758), .B2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n292), .B1(new_n753), .B2(new_n831), .C1(new_n402), .C2(new_n777), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n228), .B2(new_n774), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n999), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n795), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n963), .A2(new_n798), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n803), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n799), .B1(new_n211), .B2(new_n466), .C1(new_n1012), .C2(new_n244), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n820), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n990), .A2(new_n1014), .ZN(G387));
  OR2_X1    g0815(.A1(new_n985), .A2(new_n745), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n700), .A3(new_n986), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n765), .A2(new_n466), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n374), .B(new_n1018), .C1(G68), .C2(new_n761), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n774), .A2(new_n220), .B1(new_n753), .B2(new_n832), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n229), .B2(new_n789), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n779), .A2(G50), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G159), .A2(new_n770), .B1(new_n757), .B2(new_n261), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G311), .A2(new_n757), .B1(new_n770), .B2(G322), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n589), .B2(new_n762), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G317), .B2(new_n779), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT48), .Z(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n998), .B2(new_n765), .C1(new_n766), .C2(new_n777), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT49), .Z(new_n1030));
  INV_X1    g0830(.A(G326), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n374), .B1(new_n753), .B2(new_n1031), .C1(new_n579), .C2(new_n774), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n795), .ZN(new_n1034));
  AOI21_X1  g0834(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n470), .A2(new_n279), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n702), .B(new_n1035), .C1(new_n1036), .C2(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT50), .B2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n803), .B1(new_n241), .B2(new_n502), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n702), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n801), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n211), .A2(G107), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n799), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n692), .A2(new_n808), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1034), .A2(new_n820), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT113), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n985), .A2(new_n989), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1017), .A2(new_n1047), .A3(new_n1048), .ZN(G393));
  AOI22_X1  g0849(.A1(G107), .A2(new_n775), .B1(new_n754), .B2(G322), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n758), .B2(new_n589), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G311), .A2(new_n779), .B1(new_n770), .B2(G317), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  AOI21_X1  g0853(.A(new_n292), .B1(new_n791), .B2(G116), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n766), .C2(new_n762), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1051), .B(new_n1055), .C1(G283), .C2(new_n789), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n374), .B1(new_n791), .B2(G77), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G150), .A2(new_n770), .B1(new_n779), .B2(G159), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1057), .B1(new_n217), .B2(new_n777), .C1(new_n1058), .C2(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n757), .A2(G50), .B1(G87), .B2(new_n775), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n471), .C2(new_n762), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1059), .B(new_n1062), .C1(G143), .C2(new_n754), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n795), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n799), .B1(new_n220), .B2(new_n211), .C1(new_n1012), .C2(new_n248), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n820), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n798), .C2(new_n973), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n701), .B1(new_n980), .B2(new_n986), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n987), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n980), .B1(G1), .B2(new_n748), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(G390));
  NAND3_X1  g0874(.A1(new_n939), .A2(new_n670), .A3(new_n853), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n852), .A2(G330), .A3(new_n814), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n895), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n744), .A2(new_n818), .A3(new_n895), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n717), .A2(new_n688), .A3(new_n814), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n923), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n895), .B1(new_n744), .B2(new_n818), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n852), .A2(new_n915), .A3(G330), .A4(new_n814), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n922), .A2(new_n923), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1075), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n932), .B(new_n934), .C1(new_n930), .C2(new_n924), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1080), .A2(new_n915), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n889), .A3(new_n931), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1091), .A3(new_n1078), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1088), .B(new_n1092), .C1(new_n1093), .C2(new_n1084), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n700), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1075), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1089), .A2(new_n1078), .A3(new_n1091), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1094), .A2(KEYINPUT115), .A3(new_n700), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1097), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n932), .A2(new_n934), .A3(new_n796), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT54), .B(G143), .Z(new_n1107));
  AOI22_X1  g0907(.A1(G132), .A2(new_n779), .B1(new_n761), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n786), .C1(new_n1003), .C2(new_n765), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G50), .A2(new_n775), .B1(new_n754), .B2(G125), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n292), .B(new_n1111), .C1(new_n758), .C2(new_n831), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n789), .A2(G150), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1110), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G97), .A2(new_n761), .B1(new_n779), .B2(G116), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n998), .B2(new_n786), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G87), .A2(new_n789), .B1(new_n754), .B2(G294), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n202), .B2(new_n765), .C1(new_n758), .C2(new_n487), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1117), .A2(new_n1119), .A3(new_n292), .A4(new_n837), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n795), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n844), .A2(new_n262), .ZN(new_n1122));
  AND4_X1   g0922(.A1(new_n820), .A2(new_n1106), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n989), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1105), .A2(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1075), .B1(new_n1124), .B2(new_n1088), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n314), .A2(new_n281), .A3(new_n860), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n281), .A2(new_n860), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n308), .A2(new_n313), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n919), .B2(G330), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n903), .B(new_n1136), .C1(new_n917), .C2(new_n918), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1129), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n936), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n902), .B2(new_n903), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n919), .A2(G330), .A3(new_n1137), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1129), .A3(new_n937), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1128), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1127), .B1(new_n1146), .B2(KEYINPUT57), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n937), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1143), .A3(new_n936), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1148), .A2(new_n1149), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n701), .B1(new_n1150), .B2(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n937), .B1(new_n1144), .B2(new_n1129), .ZN(new_n1153));
  AOI211_X1 g0953(.A(KEYINPUT116), .B(new_n936), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(KEYINPUT117), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1147), .A2(new_n1151), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1136), .A2(new_n796), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n279), .B1(new_n372), .B2(G41), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1107), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n762), .A2(new_n831), .B1(new_n777), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G125), .A2(new_n770), .B1(new_n779), .B2(G128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n835), .B2(new_n758), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G150), .C2(new_n791), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT59), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G33), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n754), .B2(G124), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n1003), .C2(new_n774), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1160), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1002), .B1(new_n762), .B2(new_n466), .C1(new_n579), .C2(new_n786), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n774), .A2(new_n402), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n785), .A2(new_n487), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n777), .A2(new_n228), .B1(new_n753), .B2(new_n998), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n757), .A2(G97), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1176), .A2(new_n288), .A3(new_n374), .A4(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT58), .Z(new_n1179));
  OAI21_X1  g0979(.A(new_n795), .B1(new_n1171), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n844), .A2(new_n279), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1159), .A2(new_n820), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n989), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1158), .A2(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n895), .A2(new_n796), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1173), .A2(new_n374), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT118), .Z(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n832), .B2(new_n762), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n770), .A2(G132), .B1(G159), .B2(new_n789), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n279), .B2(new_n765), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n785), .A2(new_n831), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n758), .A2(new_n1161), .B1(new_n1109), .B2(new_n753), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1018), .B1(new_n757), .B2(G116), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G97), .A2(new_n789), .B1(new_n754), .B2(G303), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n374), .A3(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G107), .A2(new_n761), .B1(new_n779), .B2(G283), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n766), .B2(new_n786), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G77), .C2(new_n775), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n795), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n844), .A2(new_n217), .ZN(new_n1203));
  AND4_X1   g1003(.A1(new_n820), .A2(new_n1187), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1098), .B2(new_n989), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(new_n972), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1207), .B2(new_n1088), .ZN(G381));
  INV_X1    g1008(.A(KEYINPUT119), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1105), .B2(new_n1125), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1105), .A2(new_n1209), .A3(new_n1125), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G375), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(G381), .A2(G384), .ZN(new_n1215));
  INV_X1    g1015(.A(G390), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n990), .A3(new_n1014), .ZN(new_n1217));
  OR2_X1    g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1214), .A2(new_n1215), .A3(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n1214), .A2(new_n677), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT120), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(G409));
  NAND2_X1  g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1218), .A2(KEYINPUT124), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT124), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT125), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1228), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT125), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1226), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G387), .A2(G390), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1229), .A2(new_n1232), .A3(new_n1217), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(G390), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G387), .A2(new_n1235), .A3(new_n1216), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n1228), .C2(new_n1227), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1158), .A2(G378), .A3(new_n1185), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n989), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1182), .B(new_n1244), .C1(new_n1155), .C2(new_n972), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1212), .B2(new_n1210), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n677), .A2(G213), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1206), .A2(KEYINPUT60), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1082), .A2(new_n1087), .A3(new_n1075), .A4(KEYINPUT60), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1100), .A2(new_n700), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1205), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G384), .B(new_n1205), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n677), .A2(KEYINPUT122), .A3(G213), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT123), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1255), .A2(new_n1260), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1262), .B(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1249), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1247), .A2(new_n1267), .A3(new_n1248), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT121), .B1(new_n1269), .B2(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1247), .A2(KEYINPUT121), .A3(new_n1267), .A4(new_n1248), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1241), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT121), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(KEYINPUT63), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1268), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(new_n1278), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1279), .A2(new_n1265), .A3(new_n1240), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(G405));
  OAI21_X1  g1082(.A(G375), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1242), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1267), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1266), .A3(new_n1242), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1241), .B(new_n1287), .ZN(G402));
endmodule


