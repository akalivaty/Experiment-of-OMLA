//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(G8gat), .Z(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n207), .A2(KEYINPUT90), .A3(KEYINPUT15), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT90), .B1(new_n207), .B2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT92), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n213), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n216));
  OR3_X1    g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n212), .B(new_n216), .C1(new_n219), .C2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n217), .A2(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n223), .B2(new_n226), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n206), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n206), .B1(new_n223), .B2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(new_n226), .ZN(new_n235));
  INV_X1    g034(.A(new_n206), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n233), .B(KEYINPUT13), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n227), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n231), .B1(new_n242), .B2(new_n206), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n233), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT11), .B(G169gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n240), .B(new_n246), .C1(KEYINPUT93), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n234), .A2(KEYINPUT93), .A3(new_n239), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT18), .B1(new_n243), .B2(new_n233), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G148gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT77), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G148gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(G141gat), .ZN(new_n263));
  INV_X1    g062(.A(G141gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G148gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  INV_X1    g066(.A(G155gat), .ZN(new_n268));
  INV_X1    g067(.A(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n267), .B1(new_n270), .B2(KEYINPUT2), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n270), .A2(new_n267), .ZN(new_n273));
  XNOR2_X1  g072(.A(G141gat), .B(G148gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(KEYINPUT76), .C1(KEYINPUT2), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n259), .A2(G141gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT2), .B1(new_n265), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n267), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n272), .A2(new_n275), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285));
  INV_X1    g084(.A(G127gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G134gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G127gat), .ZN(new_n289));
  OAI22_X1  g088(.A1(new_n285), .A2(KEYINPUT1), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G120gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n284), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n290), .A2(new_n298), .A3(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n272), .A2(new_n275), .A3(new_n280), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT4), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n290), .A2(new_n298), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n308), .A2(new_n275), .A3(new_n272), .A4(new_n280), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n300), .A2(new_n306), .A3(new_n307), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n281), .A2(new_n299), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n309), .A3(KEYINPUT78), .ZN(new_n314));
  INV_X1    g113(.A(new_n307), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n281), .A2(new_n316), .A3(new_n299), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(new_n318), .A3(KEYINPUT5), .ZN(new_n319));
  INV_X1    g118(.A(new_n304), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n310), .B1(new_n320), .B2(new_n281), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n308), .B1(new_n281), .B2(KEYINPUT3), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n322), .B2(new_n284), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n305), .A2(KEYINPUT4), .A3(new_n308), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n321), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT0), .ZN(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT84), .A3(new_n326), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n333), .A3(new_n326), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343));
  INV_X1    g142(.A(G211gat), .ZN(new_n344));
  INV_X1    g143(.A(G218gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(KEYINPUT26), .ZN(new_n351));
  INV_X1    g150(.A(G169gat), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n350), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n358));
  INV_X1    g157(.A(G183gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT27), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(KEYINPUT27), .ZN(new_n363));
  NOR2_X1   g162(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n360), .A2(new_n362), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n359), .A2(KEYINPUT27), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n361), .A2(G183gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(G183gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n363), .A3(KEYINPUT67), .ZN(new_n371));
  AOI21_X1  g170(.A(G190gat), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n365), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT68), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G190gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n370), .A2(new_n363), .A3(KEYINPUT67), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT67), .B1(new_n370), .B2(new_n363), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT28), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(KEYINPUT68), .A3(new_n365), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n357), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(new_n352), .A3(new_n353), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT64), .B(new_n385), .C1(new_n354), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n388));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT24), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n359), .A2(new_n377), .ZN(new_n392));
  NAND3_X1  g191(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT64), .A4(new_n393), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n387), .A2(new_n388), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n388), .B1(new_n387), .B2(new_n394), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT65), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n394), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT25), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT65), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n388), .A3(new_n394), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G226gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n383), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n406), .A2(KEYINPUT29), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n357), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT68), .B1(new_n381), .B2(new_n365), .ZN(new_n412));
  INV_X1    g211(.A(new_n365), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n375), .B(new_n413), .C1(new_n380), .C2(KEYINPUT28), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n395), .A2(new_n396), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n349), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n409), .B1(new_n383), .B2(new_n403), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n415), .A2(new_n406), .A3(new_n416), .ZN(new_n422));
  INV_X1    g221(.A(new_n349), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT73), .B(new_n349), .C1(new_n408), .C2(new_n417), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND4_X1  g227(.A1(new_n420), .A2(new_n424), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n327), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT86), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n327), .A2(new_n432), .A3(KEYINPUT6), .A4(new_n334), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n341), .A2(new_n429), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n421), .A2(new_n422), .A3(new_n349), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n397), .A2(new_n402), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n415), .A2(new_n406), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n416), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n409), .B1(new_n383), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n423), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT38), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n420), .A2(new_n444), .A3(new_n424), .A4(new_n425), .ZN(new_n445));
  INV_X1    g244(.A(new_n428), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT87), .B1(new_n434), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n424), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT73), .B1(new_n441), .B2(new_n349), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT74), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n420), .A2(new_n452), .A3(new_n424), .A4(new_n425), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n451), .A2(KEYINPUT37), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(new_n446), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT38), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n433), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n333), .B1(new_n327), .B2(new_n328), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n339), .B1(new_n458), .B2(new_n335), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n429), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466));
  INV_X1    g265(.A(G50gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G228gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n349), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT3), .B1(new_n473), .B2(KEYINPUT80), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT80), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n349), .A2(new_n475), .A3(new_n472), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n305), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n349), .B1(new_n284), .B2(new_n472), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n281), .A2(new_n349), .A3(new_n472), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n471), .B1(new_n281), .B2(KEYINPUT3), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n480), .A2(KEYINPUT81), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n481), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n484), .B1(new_n485), .B2(new_n478), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G22gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n479), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n479), .B2(new_n487), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n465), .B(new_n470), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n491), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n489), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n470), .B1(new_n495), .B2(new_n465), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(KEYINPUT82), .A3(new_n489), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n451), .A2(new_n453), .A3(new_n446), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n449), .A2(new_n450), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n428), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n429), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n321), .A2(new_n300), .A3(new_n325), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n315), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n314), .A2(new_n317), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n307), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(KEYINPUT39), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT39), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n510), .A3(new_n315), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n509), .A2(KEYINPUT40), .A3(new_n333), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n336), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT40), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n506), .A2(KEYINPUT39), .A3(new_n508), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n333), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n513), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT85), .B1(new_n504), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n504), .A2(new_n521), .A3(KEYINPUT85), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n464), .B(new_n498), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n496), .A2(new_n497), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n492), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n499), .A2(KEYINPUT75), .A3(new_n501), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n327), .A2(new_n334), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n340), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n529), .A2(new_n430), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n531), .A3(new_n503), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT75), .B1(new_n499), .B2(new_n501), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n304), .B1(new_n383), .B2(new_n403), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n415), .A2(new_n320), .A3(new_n437), .ZN(new_n537));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G43gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G71gat), .B(G99gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n540), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(new_n544), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n543), .B1(new_n540), .B2(KEYINPUT32), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n548), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT34), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n383), .A2(new_n403), .A3(new_n304), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n320), .B1(new_n415), .B2(new_n437), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n553), .B(new_n538), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT71), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n536), .A2(new_n537), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n538), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT34), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT71), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n558), .A2(new_n561), .A3(new_n553), .A4(new_n538), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n535), .B1(new_n552), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n551), .A2(new_n550), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n535), .A3(new_n568), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n552), .A2(new_n563), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(KEYINPUT36), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n524), .A2(new_n534), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n578));
  NOR3_X1   g377(.A1(new_n526), .A2(new_n460), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n504), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n498), .A2(new_n574), .A3(new_n569), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n583), .A2(new_n532), .A3(new_n533), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n258), .B1(new_n577), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT7), .ZN(new_n589));
  AND2_X1   g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(KEYINPUT7), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n591), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT102), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT103), .B(G85gat), .Z(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n596), .A2(new_n597), .B1(KEYINPUT8), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n603), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n242), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n235), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT41), .ZN(new_n609));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT99), .Z(new_n611));
  OAI211_X1 g410(.A(new_n606), .B(new_n608), .C1(new_n609), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n609), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n619), .A3(new_n615), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G64gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(G57gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(G57gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G71gat), .ZN(new_n632));
  INV_X1    g431(.A(G78gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n631), .A2(new_n635), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n630), .B1(KEYINPUT96), .B2(new_n628), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(KEYINPUT96), .B2(new_n628), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n642), .B(new_n626), .C1(new_n634), .C2(new_n636), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n236), .B1(new_n647), .B2(KEYINPUT21), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT21), .B1(new_n640), .B2(new_n643), .ZN(new_n649));
  XNOR2_X1  g448(.A(G127gat), .B(G155gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n648), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT97), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n652), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n623), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n644), .B1(new_n604), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n605), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n602), .B(new_n604), .C1(new_n662), .C2(new_n644), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT10), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n646), .A2(new_n605), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n661), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n661), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n664), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n587), .A2(new_n660), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n531), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(G1gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1324gat));
  XNOR2_X1  g482(.A(KEYINPUT16), .B(G8gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT107), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n660), .A2(new_n679), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n580), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n587), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(KEYINPUT106), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n691), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT108), .B1(new_n691), .B2(KEYINPUT42), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n694), .A2(G8gat), .B1(new_n688), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(G1325gat));
  NAND2_X1  g497(.A1(new_n576), .A2(KEYINPUT109), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n573), .A2(new_n700), .A3(new_n575), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n680), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n581), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n686), .A2(G15gat), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n587), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT110), .Z(G1326gat));
  NOR2_X1   g507(.A1(new_n680), .A2(new_n498), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(new_n623), .ZN(new_n712));
  INV_X1    g511(.A(new_n659), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n713), .A3(new_n678), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n587), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n531), .A2(G29gat), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n715), .A2(KEYINPUT111), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT111), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n659), .B(KEYINPUT112), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(new_n258), .A3(new_n678), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n524), .A2(new_n699), .A3(new_n534), .A4(new_n701), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n586), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT113), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n728), .A3(new_n586), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n577), .A2(new_n586), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n623), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n724), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n531), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n738), .ZN(G1328gat));
  OAI21_X1  g538(.A(G36gat), .B1(new_n737), .B2(new_n580), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n715), .A2(G36gat), .A3(new_n580), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT114), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n742), .A2(KEYINPUT114), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n740), .B(new_n745), .C1(new_n743), .C2(new_n741), .ZN(G1329gat));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n715), .A2(G43gat), .A3(new_n704), .ZN(new_n748));
  INV_X1    g547(.A(new_n702), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n725), .A2(new_n728), .A3(new_n586), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n728), .B1(new_n725), .B2(new_n586), .ZN(new_n751));
  INV_X1    g550(.A(new_n730), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n749), .B(new_n723), .C1(new_n753), .C2(new_n734), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n748), .B1(new_n754), .B2(G43gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n747), .B1(new_n755), .B2(KEYINPUT115), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n736), .B2(new_n749), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(KEYINPUT47), .C1(new_n759), .C2(new_n748), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n756), .A2(new_n760), .ZN(G1330gat));
  AOI21_X1  g560(.A(new_n467), .B1(new_n736), .B2(new_n526), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n715), .A2(G50gat), .A3(new_n498), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n751), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n660), .A2(new_n258), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n679), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT116), .Z(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n530), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n504), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT49), .B(G64gat), .Z(new_n778));
  NOR3_X1   g577(.A1(new_n772), .A2(new_n580), .A3(new_n778), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n777), .A2(KEYINPUT117), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT117), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1333gat));
  OAI21_X1  g581(.A(G71gat), .B1(new_n772), .B2(new_n702), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n581), .A2(new_n632), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1334gat));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n498), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n633), .ZN(G1335gat));
  NAND2_X1  g588(.A1(new_n731), .A2(new_n735), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n258), .A2(new_n659), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT118), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n678), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT119), .B1(new_n794), .B2(new_n531), .ZN(new_n795));
  INV_X1    g594(.A(new_n596), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n794), .A2(KEYINPUT119), .A3(new_n531), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n726), .A2(new_n623), .A3(new_n792), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n678), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n530), .A2(new_n596), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n797), .A2(new_n798), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  AND2_X1   g604(.A1(new_n790), .A2(new_n793), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n597), .B1(new_n806), .B2(new_n504), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n504), .A2(new_n597), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G92gat), .B1(new_n794), .B2(new_n580), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n811), .B(new_n812), .C1(new_n803), .C2(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n794), .B2(new_n702), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n704), .A2(G99gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n803), .B2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n806), .B2(new_n526), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n526), .A2(new_n818), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT53), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n794), .B2(new_n498), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n823), .B(new_n824), .C1(new_n803), .C2(new_n820), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1339gat));
  NAND2_X1  g625(.A1(new_n669), .A2(KEYINPUT54), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n666), .A2(new_n668), .A3(new_n661), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT120), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n666), .A2(new_n668), .A3(new_n661), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n830), .A2(new_n669), .A3(new_n831), .A4(KEYINPUT54), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n661), .C1(new_n666), .C2(new_n668), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n675), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n829), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n253), .A2(new_n257), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n832), .A4(new_n835), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n676), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n240), .A2(new_n246), .A3(new_n252), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n243), .A2(new_n233), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n237), .A2(new_n238), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n250), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n678), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n623), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n840), .A2(new_n676), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n846), .A2(new_n621), .A3(new_n622), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(new_n838), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT121), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n850), .A3(new_n838), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n258), .B1(new_n836), .B2(new_n837), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n855), .A2(new_n849), .B1(new_n678), .B2(new_n846), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n853), .B(new_n854), .C1(new_n856), .C2(new_n623), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n857), .A3(new_n721), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n769), .A2(new_n678), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n531), .A2(new_n504), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n704), .A2(new_n526), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n293), .A3(new_n258), .ZN(new_n865));
  INV_X1    g664(.A(new_n862), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n583), .B(new_n866), .C1(new_n858), .C2(new_n860), .ZN(new_n867));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n839), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n865), .A2(new_n868), .ZN(G1340gat));
  NOR3_X1   g668(.A1(new_n864), .A2(new_n291), .A3(new_n679), .ZN(new_n870));
  AOI21_X1  g669(.A(G120gat), .B1(new_n867), .B2(new_n678), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n864), .B2(new_n721), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n867), .A2(new_n286), .A3(new_n713), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1342gat));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n712), .A2(G134gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n867), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n867), .A2(new_n877), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n864), .B2(new_n712), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n880), .A2(new_n881), .A3(new_n883), .A4(new_n884), .ZN(G1343gat));
  XOR2_X1   g684(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n749), .A2(new_n866), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n498), .B1(new_n858), .B2(new_n860), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n854), .B1(new_n856), .B2(new_n623), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n859), .B1(new_n891), .B2(new_n659), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n498), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n839), .B(new_n888), .C1(new_n890), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n866), .B1(new_n858), .B2(new_n860), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n749), .A2(new_n498), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n258), .A2(G141gat), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n887), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n886), .B(new_n900), .C1(new_n895), .C2(G141gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1344gat));
  NAND2_X1  g703(.A1(new_n897), .A2(new_n898), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT59), .B1(new_n905), .B2(new_n679), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n260), .A3(new_n262), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n679), .A2(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n888), .B(new_n908), .C1(new_n890), .C2(new_n894), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n526), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n659), .B1(new_n848), .B2(new_n851), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n498), .B1(new_n860), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(KEYINPUT57), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT124), .B(new_n893), .C1(new_n892), .C2(new_n498), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(new_n678), .A3(new_n888), .ZN(new_n917));
  NAND2_X1  g716(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n907), .B(new_n909), .C1(new_n917), .C2(new_n918), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n890), .A2(new_n894), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(new_n749), .A3(new_n866), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n721), .A2(new_n268), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n905), .A2(KEYINPUT125), .A3(new_n659), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(G155gat), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT125), .B1(new_n905), .B2(new_n659), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n921), .A2(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1346gat));
  INV_X1    g725(.A(new_n905), .ZN(new_n927));
  AOI21_X1  g726(.A(G162gat), .B1(new_n927), .B2(new_n623), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n712), .A2(new_n269), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n921), .B2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n580), .A2(new_n530), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n861), .A2(new_n863), .A3(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n352), .A3(new_n258), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n861), .A2(new_n931), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n583), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n839), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n936), .B2(new_n352), .ZN(G1348gat));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n353), .A3(new_n678), .ZN(new_n938));
  OAI21_X1  g737(.A(G176gat), .B1(new_n932), .B2(new_n679), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1349gat));
  OAI211_X1 g739(.A(new_n935), .B(new_n713), .C1(new_n378), .C2(new_n379), .ZN(new_n941));
  OAI21_X1  g740(.A(G183gat), .B1(new_n932), .B2(new_n721), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT60), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n945), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n377), .A3(new_n623), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n861), .A2(new_n623), .A3(new_n863), .A4(new_n931), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G190gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n953), .A3(G190gat), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  AND2_X1   g756(.A1(new_n702), .A2(new_n931), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n889), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n839), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n916), .A2(new_n839), .A3(new_n958), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n960), .B2(new_n963), .ZN(G1352gat));
  INV_X1    g763(.A(G204gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n959), .A2(new_n965), .A3(new_n678), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n916), .A2(new_n678), .A3(new_n958), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n967), .B(new_n968), .C1(new_n965), .C2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n344), .A3(new_n713), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n916), .A2(new_n713), .A3(new_n958), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n345), .A3(new_n623), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n916), .A2(new_n623), .A3(new_n958), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n345), .ZN(G1355gat));
endmodule


