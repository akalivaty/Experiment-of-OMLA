//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n202), .A2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208));
  OAI21_X1  g007(.A(G8gat), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n206), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n211), .A2(new_n216), .A3(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(G36gat), .B1(new_n213), .B2(new_n214), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT15), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  INV_X1    g025(.A(new_n224), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(KEYINPUT15), .C1(new_n222), .C2(new_n219), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n226), .B1(new_n225), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n210), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n232), .B(KEYINPUT88), .Z(new_n233));
  OAI211_X1 g032(.A(new_n206), .B(G8gat), .C1(new_n208), .C2(new_n207), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n209), .A2(new_n203), .A3(new_n205), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(new_n228), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT11), .B(G169gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n233), .A4(new_n238), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n233), .B(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n235), .A3(new_n225), .A4(new_n228), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n238), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n241), .A2(new_n246), .A3(new_n247), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT90), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n239), .B2(new_n240), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT90), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n246), .A4(new_n247), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n246), .B1(new_n255), .B2(new_n247), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT39), .ZN(new_n263));
  INV_X1    g062(.A(G155gat), .ZN(new_n264));
  INV_X1    g063(.A(G162gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT2), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G155gat), .B(G162gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G141gat), .B(G148gat), .Z(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n266), .C1(new_n272), .C2(new_n270), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(KEYINPUT1), .B2(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n274), .A2(new_n281), .A3(new_n276), .A4(new_n283), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n263), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n286), .B(KEYINPUT4), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT74), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n277), .A2(KEYINPUT3), .B1(new_n281), .B2(new_n283), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(KEYINPUT75), .A3(new_n298), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n291), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n289), .B1(new_n303), .B2(new_n288), .ZN(new_n304));
  XOR2_X1   g103(.A(G1gat), .B(G29gat), .Z(new_n305));
  XNOR2_X1  g104(.A(G57gat), .B(G85gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  AND3_X1   g108(.A1(new_n297), .A2(KEYINPUT75), .A3(new_n298), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT75), .B1(new_n297), .B2(new_n298), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n290), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n288), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n263), .A3(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n304), .A2(KEYINPUT40), .A3(new_n309), .A4(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n309), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT77), .B(KEYINPUT5), .C1(new_n287), .C2(new_n288), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n288), .B1(new_n285), .B2(new_n286), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT5), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n301), .A2(new_n302), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n286), .B2(KEYINPUT4), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n286), .A2(KEYINPUT4), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n286), .A2(new_n324), .A3(KEYINPUT4), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n313), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n322), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n313), .A2(KEYINPUT5), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n290), .B(new_n331), .C1(new_n310), .C2(new_n311), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n316), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n315), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT64), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT24), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(G183gat), .A3(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT23), .ZN(new_n348));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(G169gat), .B2(G176gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  INV_X1    g154(.A(new_n339), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n345), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n352), .A2(new_n355), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n354), .A2(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(G183gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT65), .A3(KEYINPUT27), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(G183gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n368), .A2(new_n369), .B1(new_n370), .B2(new_n347), .ZN(new_n371));
  NOR4_X1   g170(.A1(KEYINPUT67), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n341), .B(new_n367), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(KEYINPUT27), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n365), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n365), .A3(KEYINPUT66), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n373), .B1(new_n381), .B2(KEYINPUT28), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n338), .B1(new_n359), .B2(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n371), .A2(new_n372), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n367), .A2(new_n341), .ZN(new_n385));
  AOI21_X1  g184(.A(G190gat), .B1(new_n377), .B2(new_n378), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT28), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n353), .A2(new_n357), .A3(KEYINPUT25), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n352), .B1(new_n340), .B2(new_n345), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(KEYINPUT25), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n383), .B1(new_n392), .B2(new_n338), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT22), .ZN(new_n394));
  INV_X1    g193(.A(G211gat), .ZN(new_n395));
  INV_X1    g194(.A(G218gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT70), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT70), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  XNOR2_X1  g199(.A(G197gat), .B(G204gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(G211gat), .B(G218gat), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n402), .B(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n336), .B1(new_n393), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n337), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n402), .B(new_n403), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n337), .B1(new_n388), .B2(new_n391), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT72), .B(new_n337), .C1(new_n388), .C2(new_n391), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n410), .B(new_n411), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n393), .A2(new_n336), .A3(new_n405), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n427), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n304), .A2(new_n309), .A3(new_n314), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT40), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n335), .A2(new_n426), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n297), .A2(new_n408), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n405), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT29), .B1(new_n295), .B2(new_n296), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT81), .B1(new_n437), .B2(new_n411), .ZN(new_n438));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n292), .B1(new_n405), .B2(KEYINPUT29), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n277), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n436), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n439), .B(KEYINPUT80), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n437), .A2(new_n411), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n411), .A2(new_n408), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n445), .A2(new_n292), .B1(new_n276), .B2(new_n274), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n433), .B1(new_n448), .B2(G22gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(G78gat), .B(G106gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G22gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n442), .B2(new_n447), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n442), .A2(new_n454), .A3(new_n447), .ZN(new_n456));
  OAI22_X1  g255(.A1(new_n449), .A2(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n455), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n447), .A3(new_n454), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n433), .A3(new_n459), .A4(new_n452), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n424), .A2(KEYINPUT37), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n425), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n410), .A2(new_n411), .A3(new_n383), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n383), .A2(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n412), .A2(new_n413), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n466), .A2(new_n467), .B1(new_n337), .B2(new_n409), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT83), .B(new_n465), .C1(new_n468), .C2(new_n411), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n393), .A2(new_n405), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT38), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n329), .B1(new_n311), .B2(new_n310), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n317), .A2(new_n321), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n332), .A3(new_n309), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n334), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n316), .B(new_n480), .C1(new_n330), .C2(new_n333), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n475), .A2(new_n482), .A3(new_n483), .A4(new_n423), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n417), .A2(KEYINPUT37), .A3(new_n418), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n464), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n432), .B(new_n462), .C1(new_n484), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n482), .A2(new_n483), .ZN(new_n490));
  INV_X1    g289(.A(new_n487), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n464), .A2(new_n474), .B1(new_n419), .B2(new_n422), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n432), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n407), .A2(new_n284), .ZN(new_n497));
  NAND2_X1  g296(.A1(G227gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n284), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n388), .A2(new_n391), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT34), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n497), .A2(new_n503), .A3(new_n498), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n500), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n388), .B2(new_n391), .ZN(new_n507));
  OAI211_X1 g306(.A(G227gat), .B(G233gat), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G15gat), .B(G43gat), .Z(new_n511));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n505), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n498), .B1(new_n497), .B2(new_n500), .ZN(new_n515));
  INV_X1    g314(.A(new_n509), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n502), .A3(new_n504), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(KEYINPUT32), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n514), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n514), .B2(new_n518), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n426), .A2(new_n428), .B1(new_n482), .B2(new_n483), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n529), .B(new_n530), .C1(new_n462), .C2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n496), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n518), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n519), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n518), .A3(new_n520), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n457), .A2(new_n460), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT86), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT86), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n523), .A2(new_n540), .A3(new_n460), .A4(new_n457), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n543));
  INV_X1    g342(.A(new_n538), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n531), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT85), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(new_n531), .A3(new_n548), .A4(new_n545), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n543), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n262), .B1(new_n534), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G57gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(G64gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(KEYINPUT94), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(KEYINPUT94), .B2(new_n554), .ZN(new_n556));
  INV_X1    g355(.A(G71gat), .ZN(new_n557));
  INV_X1    g356(.A(G78gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT9), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT92), .B1(new_n563), .B2(new_n553), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(G57gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n554), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  OR3_X1    g368(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n570), .A2(new_n571), .B1(G71gat), .B2(G78gat), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n568), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n561), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT96), .ZN(new_n579));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n236), .B1(new_n576), .B2(KEYINPUT21), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n585), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n584), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT101), .B(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n591), .A2(new_n592), .B1(KEYINPUT8), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  OR2_X1    g396(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n601));
  AND2_X1   g400(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n602));
  NOR2_X1   g401(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n594), .A2(new_n596), .A3(new_n600), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n604), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT101), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G85gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n610), .A3(new_n592), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n593), .A2(KEYINPUT8), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n595), .B1(new_n606), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n229), .B2(new_n230), .ZN(new_n616));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n605), .A2(new_n614), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(new_n237), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT102), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n622), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n617), .A2(new_n618), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  XOR2_X1   g427(.A(G134gat), .B(G162gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n626), .A2(new_n630), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n575), .A2(new_n615), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  XNOR2_X1  g441(.A(G57gat), .B(G64gat), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT9), .B1(new_n643), .B2(new_n566), .ZN(new_n644));
  INV_X1    g443(.A(new_n567), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n572), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT93), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n561), .A3(new_n620), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n642), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n649), .A2(new_n620), .A3(KEYINPUT10), .A4(new_n561), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n640), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT103), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n639), .B1(new_n641), .B2(new_n650), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n638), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n653), .A2(new_n655), .A3(new_n638), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n590), .A2(new_n634), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n551), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n490), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(G1gat), .Z(G1324gat));
  INV_X1    g463(.A(new_n426), .ZN(new_n665));
  INV_X1    g464(.A(new_n428), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(G8gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n669), .ZN(new_n673));
  MUX2_X1   g472(.A(new_n671), .B(new_n673), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g473(.A1(new_n529), .A2(new_n530), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n661), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n524), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n661), .B2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n462), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  XOR2_X1   g481(.A(new_n584), .B(new_n589), .Z(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n659), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT105), .B1(new_n258), .B2(new_n260), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686));
  AOI211_X1 g485(.A(new_n686), .B(new_n259), .C1(new_n254), .C2(new_n257), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n633), .B1(new_n534), .B2(new_n550), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT106), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n543), .A2(new_n547), .A3(new_n549), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n532), .B1(new_n489), .B2(new_n495), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n634), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n691), .B(new_n634), .C1(new_n693), .C2(new_n694), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n534), .A2(new_n550), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n691), .A4(new_n634), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n689), .B1(new_n698), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n662), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n551), .A2(new_n634), .A3(new_n684), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(G29gat), .A3(new_n662), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n706), .B2(new_n668), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n708), .A2(G36gat), .A3(new_n668), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1329gat));
  NOR3_X1   g515(.A1(new_n708), .A2(G43gat), .A3(new_n524), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n676), .B(new_n689), .C1(new_n698), .C2(new_n704), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  OAI21_X1  g520(.A(G43gat), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n705), .A2(new_n721), .A3(new_n675), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n718), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n705), .A2(new_n461), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G50gat), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n462), .A2(G50gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n708), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n729), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  AOI211_X1 g534(.A(KEYINPUT48), .B(new_n733), .C1(new_n730), .C2(G50gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  XOR2_X1   g536(.A(new_n490), .B(KEYINPUT109), .Z(new_n738));
  INV_X1    g537(.A(new_n659), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n590), .A2(new_n634), .A3(new_n739), .A4(new_n688), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n701), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g541(.A1(new_n701), .A2(new_n740), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT110), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n667), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT49), .B(G64gat), .Z(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(G1333gat));
  NAND3_X1  g547(.A1(new_n744), .A2(G71gat), .A3(new_n675), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n557), .B1(new_n743), .B2(new_n524), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n744), .A2(new_n461), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n683), .A2(new_n688), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n659), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n698), .B2(new_n704), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n490), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n755), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT51), .B1(new_n690), .B2(new_n755), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n659), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n490), .A2(new_n591), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n758), .A2(new_n591), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  NAND4_X1  g563(.A1(new_n761), .A2(new_n592), .A3(new_n667), .A4(new_n659), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n668), .B(new_n756), .C1(new_n698), .C2(new_n704), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n592), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n766), .B2(new_n592), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n769), .A3(KEYINPUT52), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  OAI221_X1 g570(.A(new_n765), .B1(new_n768), .B2(new_n771), .C1(new_n766), .C2(new_n592), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n761), .A2(new_n523), .A3(new_n659), .ZN(new_n774));
  INV_X1    g573(.A(G99gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n676), .A2(new_n775), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n774), .A2(new_n775), .B1(new_n757), .B2(new_n776), .ZN(G1338gat));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(KEYINPUT53), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n757), .A2(new_n461), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G106gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n739), .A2(new_n462), .A3(G106gat), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT112), .Z(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n759), .B2(new_n760), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n778), .A2(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n780), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n779), .B(new_n787), .C1(new_n781), .C2(G106gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(G1339gat));
  NAND2_X1  g590(.A1(new_n651), .A2(new_n652), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n639), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT103), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT103), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n653), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n638), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n641), .A2(new_n642), .A3(new_n650), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n652), .A2(new_n640), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT54), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n802), .A2(KEYINPUT114), .A3(new_n653), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n652), .A2(new_n640), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n795), .B1(new_n805), .B2(new_n651), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT55), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n658), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n658), .C1(new_n799), .C2(new_n808), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n803), .A2(new_n807), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n799), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n810), .A2(new_n688), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n238), .A2(new_n250), .A3(new_n249), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n231), .A2(new_n238), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n233), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n254), .A2(new_n257), .B1(new_n819), .B2(new_n245), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n659), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n634), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n637), .B1(new_n654), .B2(new_n795), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT114), .B1(new_n802), .B2(new_n653), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n793), .A2(new_n806), .A3(new_n804), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n813), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n657), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n815), .B1(new_n827), .B2(new_n811), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n819), .A2(new_n245), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n258), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n820), .A2(KEYINPUT116), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n634), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n812), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n828), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n590), .B1(new_n822), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n688), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n683), .A2(new_n633), .A3(new_n739), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n461), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(new_n490), .A3(new_n668), .A4(new_n523), .ZN(new_n841));
  INV_X1    g640(.A(G113gat), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(new_n262), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n839), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n738), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n539), .A2(new_n541), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n668), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n688), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n843), .B1(new_n849), .B2(new_n842), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n841), .A2(new_n851), .A3(new_n739), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n659), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n855), .A3(new_n683), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n841), .B2(new_n590), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  INV_X1    g657(.A(G134gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n667), .A2(new_n633), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT117), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n847), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n841), .B2(new_n633), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n675), .A2(new_n662), .A3(new_n667), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n462), .B1(new_n837), .B2(new_n839), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n660), .A2(new_n838), .ZN(new_n872));
  INV_X1    g671(.A(new_n836), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n827), .A2(new_n261), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n799), .A2(new_n814), .ZN(new_n875));
  XNOR2_X1  g674(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n821), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n633), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n683), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT57), .B(new_n461), .C1(new_n872), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n870), .A2(new_n869), .A3(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n261), .B(new_n868), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n675), .A2(new_n462), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n262), .A2(G141gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n845), .A2(new_n668), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n867), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT120), .B(new_n891), .C1(new_n885), .C2(G141gat), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n688), .B(new_n868), .C1(new_n883), .C2(new_n884), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n845), .A2(new_n887), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n667), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n895), .A2(G141gat), .B1(new_n897), .B2(new_n888), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n893), .A2(new_n894), .B1(new_n890), .B2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n868), .B1(new_n883), .B2(new_n884), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n900), .B(G148gat), .C1(new_n901), .C2(new_n739), .ZN(new_n902));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n870), .A2(new_n904), .ZN(new_n905));
  NOR4_X1   g704(.A1(new_n590), .A2(new_n261), .A3(new_n634), .A4(new_n659), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(new_n461), .C1(new_n881), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n868), .A2(new_n659), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n902), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n897), .A2(new_n903), .A3(new_n659), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1345gat));
  OAI211_X1 g712(.A(new_n683), .B(new_n868), .C1(new_n883), .C2(new_n884), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G155gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n264), .A3(new_n683), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(KEYINPUT121), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n901), .B2(new_n633), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n861), .A2(new_n265), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n896), .B2(new_n923), .ZN(G1347gat));
  AOI21_X1  g723(.A(new_n490), .B1(new_n837), .B2(new_n839), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n667), .A3(new_n846), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT122), .Z(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n688), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n738), .A2(new_n668), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n524), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n840), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n261), .A2(G169gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  INV_X1    g732(.A(G176gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n927), .A2(new_n934), .A3(new_n659), .ZN(new_n935));
  INV_X1    g734(.A(new_n931), .ZN(new_n936));
  OAI21_X1  g735(.A(G176gat), .B1(new_n936), .B2(new_n739), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1349gat));
  AOI21_X1  g737(.A(new_n363), .B1(new_n931), .B2(new_n683), .ZN(new_n939));
  INV_X1    g738(.A(new_n379), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n926), .A2(new_n940), .A3(new_n590), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g742(.A(new_n380), .B1(new_n931), .B2(new_n634), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT61), .Z(new_n945));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n380), .A3(new_n634), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n929), .A2(new_n675), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n907), .B(new_n949), .C1(new_n870), .C2(new_n904), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT124), .B1(new_n950), .B2(new_n262), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G197gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n950), .A2(KEYINPUT124), .A3(new_n262), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n925), .A2(new_n667), .A3(new_n887), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n838), .A2(G197gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT123), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n948), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n957), .B(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n961), .B(KEYINPUT125), .C1(new_n953), .C2(new_n952), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n955), .A2(new_n964), .A3(new_n659), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n950), .B2(new_n739), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n395), .A3(new_n683), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n950), .A2(new_n590), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n395), .B1(KEYINPUT126), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g774(.A1(new_n970), .A2(new_n975), .B1(new_n971), .B2(KEYINPUT63), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n969), .B1(new_n973), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n950), .B2(new_n633), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n955), .A2(new_n396), .A3(new_n634), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


