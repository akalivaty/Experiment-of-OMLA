//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G221), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(new_n187), .A3(G953), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n191), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n201));
  OR3_X1    g015(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G146), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G146), .B1(new_n201), .B2(new_n202), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(G119), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT69), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT24), .B(G110), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n204), .A2(new_n205), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT69), .B(G119), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n214), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT77), .A3(new_n206), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n210), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n218), .B1(G110), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G110), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n230), .A3(new_n227), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n216), .A2(new_n217), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n225), .A2(KEYINPUT78), .A3(new_n230), .A4(new_n227), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G125), .B(G140), .ZN(new_n237));
  INV_X1    g051(.A(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n203), .A2(new_n239), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n196), .B(new_n229), .C1(new_n236), .C2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(G128), .B1(new_n212), .B2(new_n214), .ZN(new_n242));
  AOI22_X1  g056(.A1(KEYINPUT77), .A2(new_n242), .B1(new_n215), .B2(KEYINPUT23), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n243), .A2(new_n221), .B1(KEYINPUT23), .B2(new_n226), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT78), .B1(new_n244), .B2(new_n230), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n235), .A2(new_n234), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n229), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT79), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n195), .B1(new_n241), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n248), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n194), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT25), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n256), .B(G902), .C1(new_n250), .C2(new_n252), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n190), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n188), .A2(new_n254), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT80), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT2), .B(G113), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n212), .A2(new_n214), .A3(G116), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(G116), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n211), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT70), .B1(new_n220), .B2(G116), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n266), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n220), .A2(KEYINPUT70), .A3(G116), .ZN(new_n272));
  INV_X1    g086(.A(new_n264), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT71), .A2(G116), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT71), .A2(G116), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G119), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT11), .B1(new_n283), .B2(G137), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  INV_X1    g099(.A(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n286), .B2(G134), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(KEYINPUT65), .A3(G137), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G131), .ZN(new_n293));
  INV_X1    g107(.A(G131), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n288), .A2(new_n294), .A3(new_n290), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G143), .B(G146), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT64), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n238), .A2(G143), .ZN(new_n300));
  INV_X1    g114(.A(G143), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G146), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  OR2_X1    g119(.A1(KEYINPUT0), .A2(G128), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n297), .A2(KEYINPUT0), .A3(G128), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n299), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n283), .A2(G137), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n286), .A2(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT1), .B1(new_n301), .B2(G146), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n314), .A2(KEYINPUT67), .B1(new_n207), .B2(new_n209), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n300), .A2(new_n316), .A3(KEYINPUT1), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n297), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n300), .A2(new_n302), .A3(new_n319), .A4(G128), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n295), .B(new_n313), .C1(new_n318), .C2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n281), .A2(new_n282), .A3(new_n310), .A4(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G210), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT27), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n295), .A2(new_n313), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n207), .A2(new_n209), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n317), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n303), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n320), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n295), .A2(KEYINPUT66), .A3(new_n313), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n310), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n299), .A2(new_n307), .A3(new_n308), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n293), .B2(new_n295), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n321), .B1(new_n336), .B2(new_n303), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n331), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT30), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI221_X4 g161(.A(KEYINPUT73), .B1(new_n281), .B2(new_n282), .C1(new_n342), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n281), .A2(new_n282), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n330), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT31), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n328), .B(KEYINPUT74), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT75), .B1(new_n310), .B2(new_n322), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n310), .A2(KEYINPUT75), .A3(new_n322), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT28), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n340), .A2(new_n310), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(new_n323), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n356), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT31), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(new_n330), .C1(new_n348), .C2(new_n352), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G472), .A2(G902), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT32), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G472), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n372));
  INV_X1    g186(.A(new_n323), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n281), .A2(new_n282), .B1(new_n340), .B2(new_n310), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT28), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n344), .B2(new_n346), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n359), .A3(new_n281), .A4(new_n282), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n361), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n379), .A3(new_n355), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n350), .A2(new_n351), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n350), .A2(new_n349), .A3(new_n351), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n373), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n372), .B(new_n380), .C1(new_n384), .C2(new_n328), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT72), .B1(new_n270), .B2(new_n278), .ZN(new_n387));
  OAI22_X1  g201(.A1(new_n386), .A2(new_n387), .B1(new_n344), .B2(new_n346), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n323), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT28), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(KEYINPUT29), .A3(new_n379), .A4(new_n328), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(new_n254), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n371), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n370), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n369), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n367), .A2(new_n365), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n382), .A2(new_n383), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n366), .B1(new_n399), .B2(new_n330), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n263), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n403));
  NOR2_X1   g217(.A1(G475), .A2(G902), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n324), .A2(G143), .A3(G214), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G143), .B1(new_n324), .B2(G214), .ZN(new_n407));
  OAI21_X1  g221(.A(G131), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  INV_X1    g223(.A(G237), .ZN(new_n410));
  INV_X1    g224(.A(G953), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G214), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n301), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n294), .A3(new_n405), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n205), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT17), .B(G131), .C1(new_n406), .C2(new_n407), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n415), .A2(new_n203), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n405), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT18), .A2(G131), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT90), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n413), .A2(new_n423), .A3(new_n405), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n237), .A2(new_n238), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n426), .A2(new_n239), .B1(new_n419), .B2(new_n421), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G113), .B(G122), .ZN(new_n429));
  INV_X1    g243(.A(G104), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n418), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n237), .B(KEYINPUT19), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n238), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n408), .A2(new_n414), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n203), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n431), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n403), .B(new_n404), .C1(new_n432), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT20), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n418), .A2(new_n428), .A3(new_n431), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n428), .A2(new_n436), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n431), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n403), .B1(new_n442), .B2(new_n404), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n404), .B1(new_n432), .B2(new_n437), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT91), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT20), .A3(new_n438), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n416), .A2(new_n417), .A3(new_n203), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n450), .A2(new_n415), .B1(new_n425), .B2(new_n427), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT93), .B1(new_n451), .B2(new_n431), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n418), .A2(new_n428), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT93), .ZN(new_n454));
  INV_X1    g268(.A(new_n431), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n432), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n449), .B1(new_n457), .B2(G902), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT92), .B(G475), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n457), .A2(G902), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(KEYINPUT94), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n448), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n207), .A2(new_n209), .A3(G143), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n301), .A2(G128), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n283), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n466), .A2(new_n283), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G122), .ZN(new_n472));
  INV_X1    g286(.A(G122), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT95), .ZN(new_n474));
  OAI21_X1  g288(.A(G116), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G107), .ZN(new_n476));
  INV_X1    g290(.A(new_n275), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT71), .A2(G116), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(G122), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n476), .B1(new_n475), .B2(new_n479), .ZN(new_n482));
  OAI221_X1 g296(.A(new_n468), .B1(new_n469), .B2(new_n470), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n463), .A2(new_n283), .A3(new_n464), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n480), .B1(new_n484), .B2(new_n465), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n276), .B2(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT95), .B(G122), .ZN(new_n489));
  INV_X1    g303(.A(G116), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n486), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n274), .A2(new_n275), .A3(new_n473), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n487), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n475), .B(KEYINPUT96), .C1(new_n493), .C2(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT97), .B(new_n485), .C1(new_n496), .C2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n494), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n479), .A2(KEYINPUT14), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT96), .B1(new_n500), .B2(new_n475), .ZN(new_n501));
  OAI21_X1  g315(.A(G107), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n485), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n483), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT9), .B(G234), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G217), .A3(new_n411), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n483), .B(new_n508), .C1(new_n497), .C2(new_n504), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n254), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G478), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT15), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n510), .A2(KEYINPUT98), .A3(new_n254), .A4(new_n511), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT99), .A2(G952), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT99), .A2(G952), .ZN(new_n521));
  AOI21_X1  g335(.A(G953), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n187), .B2(new_n410), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n254), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT21), .B(G898), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n512), .A2(new_n516), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n462), .A2(new_n518), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G214), .B1(G237), .B2(G902), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT8), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT5), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n220), .A2(new_n534), .A3(G116), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n271), .A2(new_n272), .A3(new_n277), .ZN(new_n536));
  OAI211_X1 g350(.A(G113), .B(new_n535), .C1(new_n536), .C2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT3), .B1(new_n430), .B2(G107), .ZN(new_n538));
  AOI21_X1  g352(.A(G101), .B1(new_n430), .B2(G107), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT3), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n476), .A3(G104), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n538), .A2(new_n539), .A3(new_n541), .A4(KEYINPUT81), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n430), .B2(G107), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n430), .A2(G107), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n476), .A2(KEYINPUT82), .A3(G104), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n544), .A2(new_n545), .B1(G101), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n537), .A2(new_n278), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n537), .B2(new_n278), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n533), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n338), .A2(new_n199), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n309), .A2(G125), .ZN(new_n557));
  INV_X1    g371(.A(G224), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G953), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(KEYINPUT87), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(KEYINPUT87), .B2(new_n560), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n556), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(new_n557), .ZN(new_n564));
  INV_X1    g378(.A(new_n559), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT88), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n565), .A2(KEYINPUT88), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n564), .A2(KEYINPUT7), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n555), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n544), .A2(new_n545), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT4), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n538), .A2(new_n541), .A3(new_n548), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(G101), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n571), .A3(G101), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n386), .B2(new_n387), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n552), .A3(new_n532), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n254), .B1(new_n569), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n564), .B(new_n565), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n577), .A2(new_n552), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n532), .B(KEYINPUT86), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n578), .A2(KEYINPUT6), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G210), .B1(G237), .B2(G902), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n581), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n581), .B2(new_n587), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n531), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  XNOR2_X1  g409(.A(G110), .B(G140), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n411), .A2(G227), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n574), .A2(new_n309), .A3(new_n575), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n338), .A2(KEYINPUT10), .A3(new_n551), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n544), .A2(new_n545), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n206), .B1(new_n300), .B2(KEYINPUT1), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n320), .B1(new_n604), .B2(new_n297), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n550), .A2(G101), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n602), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n296), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n609), .A2(new_n612), .A3(new_n296), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n296), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n600), .A2(new_n601), .A3(new_n608), .A4(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n599), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n599), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n570), .A2(new_n606), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n345), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n570), .A2(new_n606), .A3(new_n605), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n296), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT12), .B1(new_n296), .B2(KEYINPUT83), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n622), .B(new_n296), .C1(KEYINPUT83), .C2(KEYINPUT12), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n618), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n595), .B(new_n254), .C1(new_n617), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n626), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n616), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n598), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT84), .B1(new_n616), .B2(new_n599), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n616), .A2(KEYINPUT84), .A3(new_n599), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n609), .A2(new_n612), .A3(new_n296), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n612), .B1(new_n609), .B2(new_n296), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n631), .B(G469), .C1(new_n632), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(G469), .A2(G902), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n628), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n192), .B1(new_n507), .B2(new_n254), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n530), .A2(new_n594), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n402), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n355), .B1(new_n375), .B2(new_n379), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n329), .B1(new_n382), .B2(new_n383), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n366), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n650), .B2(new_n354), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n651), .B2(new_n371), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n369), .B1(new_n398), .B2(new_n400), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n368), .A2(new_n254), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(KEYINPUT100), .A3(G472), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n258), .A2(new_n262), .A3(new_n641), .A4(new_n639), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n646), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n657), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n371), .B1(new_n368), .B2(new_n254), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n660), .A2(KEYINPUT100), .B1(new_n368), .B2(new_n369), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n659), .A2(KEYINPUT101), .A3(new_n652), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n439), .B(new_n446), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n451), .A2(KEYINPUT93), .A3(new_n431), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n440), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(KEYINPUT94), .A3(new_n254), .ZN(new_n667));
  INV_X1    g481(.A(new_n459), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n458), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT33), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n510), .A2(new_n671), .A3(new_n511), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n510), .A2(new_n674), .A3(new_n671), .A4(new_n511), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n508), .A2(KEYINPUT103), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n671), .B1(new_n505), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n505), .B2(new_n676), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n515), .A2(G902), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n675), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n670), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n582), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n578), .A2(KEYINPUT6), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n583), .A2(new_n584), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n588), .B1(new_n691), .B2(new_n580), .ZN(new_n692));
  INV_X1    g506(.A(new_n588), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n581), .A2(new_n587), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(new_n694), .A3(new_n528), .A4(new_n531), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n658), .A2(new_n662), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT106), .B(G104), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT105), .B(KEYINPUT34), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G6));
  AOI21_X1  g515(.A(new_n670), .B1(new_n529), .B2(new_n518), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n692), .A2(new_n531), .A3(new_n694), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .A4(new_n528), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n518), .A2(new_n529), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n462), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT107), .B1(new_n707), .B2(new_n695), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n658), .A2(new_n662), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT35), .B(G107), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G9));
  INV_X1    g526(.A(new_n642), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n706), .A2(new_n527), .A3(new_n670), .ZN(new_n714));
  INV_X1    g528(.A(new_n531), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n589), .B1(new_n691), .B2(new_n580), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(new_n591), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n241), .A2(new_n249), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n261), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n258), .A2(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n713), .A2(new_n714), .A3(new_n717), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n656), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT108), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT37), .B(G110), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G12));
  AOI21_X1  g542(.A(new_n642), .B1(new_n258), .B2(new_n721), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n653), .A2(new_n396), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n328), .B1(new_n399), .B2(new_n323), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n380), .A2(new_n372), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n392), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G472), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n401), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(G900), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n524), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n523), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n707), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n729), .A2(new_n735), .A3(new_n703), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G128), .ZN(G30));
  XOR2_X1   g555(.A(new_n738), .B(KEYINPUT39), .Z(new_n742));
  NAND2_X1  g556(.A1(new_n713), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT40), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n706), .A2(new_n670), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n722), .A2(new_n715), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n716), .A2(new_n591), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT38), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n355), .B1(new_n323), .B2(new_n388), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n254), .B1(new_n649), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G472), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n730), .A2(new_n401), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n745), .A2(new_n747), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G143), .ZN(G45));
  INV_X1    g569(.A(new_n738), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n670), .B(new_n756), .C1(new_n683), .C2(new_n684), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n735), .A3(new_n729), .A4(new_n703), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G146), .ZN(G48));
  INV_X1    g574(.A(new_n252), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n251), .A2(new_n196), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n247), .A2(KEYINPUT79), .A3(new_n248), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n761), .B1(new_n764), .B2(new_n195), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n256), .B1(new_n765), .B2(G902), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n254), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n768), .A2(new_n190), .B1(new_n261), .B2(new_n253), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n616), .B1(new_n634), .B2(new_n635), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n627), .B1(new_n770), .B2(new_n598), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n771), .B2(G902), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n628), .A3(new_n641), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n735), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n696), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT41), .B(G113), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G15));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n709), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G116), .ZN(G18));
  AND3_X1   g594(.A1(new_n735), .A2(new_n714), .A3(new_n722), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n703), .A2(new_n774), .A3(KEYINPUT109), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n692), .A2(new_n531), .A3(new_n694), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n784), .B2(new_n773), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G119), .ZN(G21));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n361), .B1(new_n323), .B2(new_n388), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n360), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n390), .A2(new_n379), .A3(KEYINPUT110), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n356), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n354), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n367), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n793), .B2(new_n354), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n369), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n660), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n798), .A2(new_n769), .A3(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n746), .A2(new_n784), .A3(new_n773), .A4(new_n527), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G122), .ZN(G24));
  AND3_X1   g617(.A1(new_n798), .A2(new_n799), .A3(new_n722), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n758), .A3(new_n786), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G125), .ZN(G27));
  NAND4_X1  g620(.A1(new_n716), .A2(new_n591), .A3(new_n641), .A4(new_n531), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n628), .A2(new_n638), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n599), .B1(new_n629), .B2(new_n616), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT112), .B1(new_n636), .B2(new_n632), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  INV_X1    g626(.A(new_n632), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n614), .A2(new_n812), .A3(new_n813), .A4(new_n633), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n595), .B(new_n810), .C1(new_n811), .C2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n808), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n810), .B1(new_n811), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(G469), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT113), .A3(new_n628), .A4(new_n638), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n807), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n401), .A2(KEYINPUT115), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n368), .A2(new_n822), .A3(new_n397), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n730), .A2(new_n821), .A3(new_n734), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n820), .A2(KEYINPUT42), .A3(new_n824), .A4(new_n769), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT116), .B1(new_n825), .B2(new_n757), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n824), .A2(new_n769), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT42), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n828), .B(new_n807), .C1(new_n816), .C2(new_n819), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n827), .A2(new_n829), .A3(new_n830), .A4(new_n758), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n758), .A2(new_n402), .A3(new_n820), .ZN(new_n832));
  XNOR2_X1  g646(.A(KEYINPUT114), .B(KEYINPUT42), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n826), .A2(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n294), .ZN(G33));
  NAND3_X1  g649(.A1(new_n402), .A2(new_n739), .A3(new_n820), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G134), .ZN(G36));
  INV_X1    g651(.A(new_n628), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n817), .A2(KEYINPUT117), .A3(KEYINPUT45), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n636), .A2(new_n632), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n810), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n839), .B(G469), .C1(KEYINPUT45), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT117), .B1(new_n817), .B2(KEYINPUT45), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n638), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT46), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n845), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n641), .ZN(new_n848));
  INV_X1    g662(.A(new_n742), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n748), .A2(new_n715), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n462), .B1(new_n683), .B2(new_n684), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT43), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(KEYINPUT118), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT118), .B(KEYINPUT43), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n656), .A2(new_n722), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT44), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(G137), .ZN(G39));
  INV_X1    g676(.A(KEYINPUT47), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n848), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n847), .A2(KEYINPUT47), .A3(new_n641), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n757), .A2(new_n851), .A3(new_n735), .A4(new_n769), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(G140), .ZN(G42));
  NAND2_X1  g683(.A1(new_n772), .A2(new_n628), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n870), .A2(KEYINPUT49), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n640), .A3(new_n715), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(KEYINPUT49), .B2(new_n870), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n753), .A2(new_n263), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OR4_X1    g689(.A1(new_n749), .A2(new_n873), .A3(new_n875), .A4(new_n853), .ZN(new_n876));
  INV_X1    g690(.A(new_n523), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n857), .A2(new_n877), .A3(new_n800), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n749), .A2(new_n531), .A3(new_n773), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(KEYINPUT50), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n807), .A2(new_n523), .A3(new_n870), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n857), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n804), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n683), .A2(new_n684), .A3(new_n670), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n885), .A3(new_n874), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n870), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n866), .B1(new_n640), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n878), .A2(new_n850), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n891), .B(KEYINPUT51), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n890), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n878), .A2(new_n786), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n874), .A2(new_n885), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n899), .B(new_n522), .C1(new_n685), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n886), .A2(new_n827), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT48), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n902), .B2(new_n904), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n901), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n895), .A2(new_n898), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n786), .A2(new_n781), .B1(new_n800), .B2(new_n801), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n748), .A2(new_n528), .A3(new_n531), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n685), .B2(new_n707), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n658), .A2(new_n662), .A3(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n723), .A2(new_n724), .B1(new_n402), .B2(new_n643), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n775), .B1(new_n696), .B2(new_n709), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n911), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n826), .A2(new_n831), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n832), .A2(new_n833), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n706), .A2(new_n670), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n756), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n851), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n922), .A3(new_n756), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n735), .A3(new_n729), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n804), .A2(new_n758), .A3(new_n820), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n836), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n918), .A2(new_n921), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n805), .A2(new_n740), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT52), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n722), .A2(new_n640), .A3(new_n738), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n816), .A2(new_n819), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n746), .A2(new_n784), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n753), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n932), .A2(new_n933), .A3(new_n759), .A4(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n759), .A2(new_n805), .A3(new_n740), .A4(new_n937), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT52), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n910), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n834), .A2(new_n917), .A3(new_n929), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n939), .B(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n805), .A2(new_n740), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT52), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n910), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT54), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT53), .A4(new_n946), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT54), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n942), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n909), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(G952), .A2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n876), .B1(new_n955), .B2(new_n956), .ZN(G75));
  NOR2_X1   g771(.A1(new_n411), .A2(G952), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT121), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n942), .A2(new_n951), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(G902), .ZN(new_n963));
  INV_X1    g777(.A(G210), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n585), .A2(new_n586), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n686), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n587), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT55), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n965), .A2(new_n970), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n960), .B1(new_n971), .B2(new_n972), .ZN(G51));
  NOR3_X1   g787(.A1(new_n963), .A2(new_n843), .A3(new_n842), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n946), .A2(KEYINPUT53), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n931), .A2(new_n941), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT53), .B1(new_n943), .B2(new_n944), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT54), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n953), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n638), .B(KEYINPUT57), .Z(new_n980));
  AOI21_X1  g794(.A(new_n771), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n974), .B1(new_n981), .B2(KEYINPUT122), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT122), .ZN(new_n983));
  INV_X1    g797(.A(new_n980), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n978), .B2(new_n953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n985), .B2(new_n771), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n958), .B1(new_n982), .B2(new_n986), .ZN(G54));
  NAND2_X1  g801(.A1(KEYINPUT58), .A2(G475), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT123), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI221_X1 g804(.A(new_n440), .B1(new_n431), .B2(new_n441), .C1(new_n963), .C2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n958), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n962), .A2(G902), .A3(new_n442), .A4(new_n989), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(G60));
  NAND3_X1  g808(.A1(new_n673), .A2(new_n675), .A3(new_n678), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT124), .ZN(new_n996));
  NAND2_X1  g810(.A1(G478), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT59), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n979), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n996), .B1(new_n954), .B2(new_n998), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n999), .A2(new_n1000), .A3(new_n960), .ZN(G63));
  NOR2_X1   g815(.A1(new_n976), .A2(new_n977), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G217), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT60), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n720), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n765), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(new_n959), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1006), .A2(KEYINPUT61), .A3(new_n959), .A4(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(G66));
  NAND2_X1  g826(.A1(new_n917), .A2(new_n411), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT125), .Z(new_n1014));
  OAI21_X1  g828(.A(G953), .B1(new_n525), .B2(new_n558), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n966), .B1(G898), .B2(new_n411), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G69));
  AOI21_X1  g832(.A(new_n411), .B1(G227), .B2(G900), .ZN(new_n1019));
  AND4_X1   g833(.A1(new_n759), .A2(new_n921), .A3(new_n836), .A4(new_n932), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n848), .A2(new_n849), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(new_n936), .A3(new_n827), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1020), .A2(new_n868), .A3(new_n861), .A4(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n350), .B(new_n433), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1023), .A2(new_n411), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n754), .A2(new_n759), .A3(new_n932), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT62), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n743), .A2(new_n851), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n402), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1029), .B1(new_n685), .B2(new_n707), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n868), .A2(new_n861), .ZN(new_n1032));
  AOI21_X1  g846(.A(G953), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1025), .B1(new_n1033), .B2(new_n1024), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1019), .B1(new_n1034), .B2(new_n736), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1035), .B1(new_n1019), .B2(new_n1034), .ZN(G72));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n1023), .B2(new_n917), .ZN(new_n1039));
  INV_X1    g853(.A(new_n328), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n384), .B(KEYINPUT127), .Z(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n949), .B(new_n1038), .C1(new_n649), .C2(new_n731), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1043), .A2(new_n992), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1031), .A2(new_n1032), .A3(new_n918), .ZN(new_n1046));
  AOI21_X1  g860(.A(KEYINPUT126), .B1(new_n1046), .B2(new_n1038), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n1047), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1046), .A2(KEYINPUT126), .A3(new_n1038), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(G57));
endmodule


