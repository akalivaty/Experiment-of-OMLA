//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1114, new_n1115;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G101), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(KEYINPUT67), .A3(G101), .A4(G2104), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n465), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n465), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT68), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(new_n485), .B2(G136), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(G162));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n478), .A2(new_n495), .A3(G138), .A4(new_n465), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(new_n505), .B(KEYINPUT71), .Z(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(G88), .B1(new_n510), .B2(G50), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT74), .B(G89), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n508), .A2(new_n518), .B1(new_n510), .B2(G51), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT73), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G168));
  NAND2_X1  g099(.A1(new_n499), .A2(new_n501), .ZN(new_n525));
  INV_X1    g100(.A(G64), .ZN(new_n526));
  INV_X1    g101(.A(G77), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n498), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(G651), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n508), .A2(G90), .B1(new_n510), .B2(G52), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  AOI22_X1  g112(.A1(new_n508), .A2(G81), .B1(new_n510), .B2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n525), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  NAND3_X1  g124(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n504), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n502), .A2(new_n507), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n551), .B(new_n553), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT78), .ZN(G299));
  XNOR2_X1  g133(.A(G168), .B(KEYINPUT79), .ZN(G286));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n554), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G87), .ZN(new_n562));
  INV_X1    g137(.A(G74), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n504), .B1(new_n525), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n510), .B2(G49), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G288));
  NAND2_X1  g141(.A1(new_n561), .A2(G86), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n525), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(G48), .A2(new_n510), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n504), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT80), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n508), .A2(G85), .B1(new_n510), .B2(G47), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(KEYINPUT80), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  INV_X1    g157(.A(G92), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n555), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n561), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n504), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n509), .B2(KEYINPUT81), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(KEYINPUT81), .B2(new_n509), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n581), .B1(new_n593), .B2(G868), .ZN(G321));
  XOR2_X1   g169(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n557), .B(KEYINPUT78), .Z(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(G868), .B2(new_n597), .ZN(G280));
  XOR2_X1   g173(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT84), .Z(G148));
  NAND2_X1  g177(.A1(new_n593), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g181(.A(new_n478), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n468), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  NOR2_X1   g186(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n612));
  AND2_X1   g187(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n615), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n616));
  INV_X1    g191(.A(G123), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n479), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n485), .B2(G135), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2096), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n614), .B(new_n620), .C1(new_n612), .C2(new_n611), .ZN(G156));
  INV_X1    g196(.A(KEYINPUT14), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT16), .B(G1341), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  AND2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  INV_X1    g221(.A(new_n638), .ZN(new_n647));
  INV_X1    g222(.A(new_n639), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(new_n642), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2096), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT20), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n660), .B(new_n662), .C1(new_n655), .C2(new_n661), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1991), .ZN(new_n666));
  INV_X1    g241(.A(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G22), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G166), .B2(new_n673), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(G1971), .ZN(new_n676));
  MUX2_X1   g251(.A(G6), .B(G305), .S(G16), .Z(new_n677));
  XOR2_X1   g252(.A(KEYINPUT32), .B(G1981), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(G16), .A2(G23), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT92), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G288), .B2(new_n673), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT33), .B(G1976), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT93), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n675), .A2(G1971), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n676), .A2(new_n679), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT34), .Z(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G25), .ZN(new_n690));
  OAI21_X1  g265(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g267(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n693));
  OAI221_X1 g268(.A(G2104), .B1(G107), .B2(new_n465), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT90), .Z(new_n695));
  INV_X1    g270(.A(G119), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n479), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n485), .A2(G131), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n690), .B1(new_n699), .B2(new_n689), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT91), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n700), .B(new_n702), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n579), .A2(new_n673), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n673), .B2(G24), .ZN(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n688), .A2(new_n703), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT36), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n673), .A2(G5), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G171), .B2(new_n673), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G1961), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT25), .ZN(new_n715));
  NAND2_X1  g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  INV_X1    g291(.A(G127), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n607), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n719));
  OAI21_X1  g294(.A(G2105), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT98), .Z(new_n722));
  AOI211_X1 g297(.A(new_n715), .B(new_n722), .C1(G139), .C2(new_n485), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(new_n689), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n689), .B2(G33), .ZN(new_n725));
  INV_X1    g300(.A(G2072), .ZN(new_n726));
  OAI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G1961), .B2(new_n712), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n713), .B(new_n727), .C1(new_n726), .C2(new_n725), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G32), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT26), .Z(new_n731));
  INV_X1    g306(.A(G105), .ZN(new_n732));
  INV_X1    g307(.A(G129), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n731), .B1(new_n732), .B2(new_n468), .C1(new_n479), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n485), .B2(G141), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT101), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n729), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n593), .A2(new_n673), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G4), .B2(new_n673), .ZN(new_n742));
  INV_X1    g317(.A(G1348), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n689), .A2(G26), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n485), .A2(G140), .ZN(new_n747));
  INV_X1    g322(.A(new_n479), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G128), .ZN(new_n749));
  OR2_X1    g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n747), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n745), .B(new_n746), .C1(new_n752), .C2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n745), .B2(new_n746), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT95), .B(G2067), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n740), .A2(new_n744), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G28), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n689), .B1(new_n759), .B2(G28), .ZN(new_n761));
  AND2_X1   g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  NOR2_X1   g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n619), .B2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(G160), .A2(G29), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G34), .Z(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(G29), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G168), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G16), .B2(G21), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n765), .B1(G2084), .B2(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n773), .B2(new_n772), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n770), .A2(G2084), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT100), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n689), .A2(G27), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G164), .B2(new_n689), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n775), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n673), .A2(G19), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n543), .B2(new_n673), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT94), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n742), .B2(new_n743), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n758), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G35), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G162), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT29), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G20), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n794), .A2(KEYINPUT23), .A3(G16), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n597), .A2(new_n673), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT23), .B1(new_n794), .B2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT102), .B(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n728), .A2(new_n788), .A3(new_n793), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n710), .A2(new_n801), .ZN(G311));
  INV_X1    g377(.A(G311), .ZN(G150));
  NAND2_X1  g378(.A1(new_n593), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT39), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n504), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT104), .B(G93), .Z(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT103), .B(G55), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n554), .A2(new_n810), .B1(new_n509), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n543), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(G860), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n814), .B2(new_n807), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT106), .ZN(new_n817));
  OAI21_X1  g392(.A(G860), .B1(new_n809), .B2(new_n812), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  NAND2_X1  g395(.A1(new_n485), .A2(G142), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT107), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n748), .A2(G130), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n465), .A2(G118), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G164), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n699), .B(new_n752), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(G162), .B(new_n619), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n610), .B(G160), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n829), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n723), .A2(new_n735), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n737), .B2(new_n723), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT108), .B(G37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n835), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g415(.A(G288), .B(G305), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G303), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n579), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT110), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT42), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(KEYINPUT42), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT109), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n593), .A2(G299), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n593), .A2(G299), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(KEYINPUT109), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT41), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n814), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n603), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n854), .A2(new_n855), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n863), .B(new_n861), .C1(new_n846), .C2(new_n847), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G868), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT111), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n813), .A2(G868), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G868), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n865), .B2(new_n866), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT111), .B1(new_n874), .B2(new_n870), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(G295));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n871), .ZN(G331));
  NAND2_X1  g452(.A1(G286), .A2(G171), .ZN(new_n878));
  NAND3_X1  g453(.A1(G301), .A2(KEYINPUT112), .A3(G168), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT112), .ZN(new_n880));
  INV_X1    g455(.A(G168), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(G171), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n883), .A2(new_n859), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n859), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n862), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n883), .B(new_n814), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n886), .B(new_n843), .C1(new_n858), .C2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT113), .ZN(new_n891));
  INV_X1    g466(.A(new_n843), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n886), .B1(new_n858), .B2(new_n887), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT43), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n884), .A2(new_n885), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(KEYINPUT41), .C1(new_n852), .C2(new_n853), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n862), .B1(new_n887), .B2(new_n849), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n843), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n837), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT44), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n894), .B2(new_n895), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(G397));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G164), .B2(G1384), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n472), .A2(new_n476), .A3(G40), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n752), .B(G2067), .Z(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(new_n735), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n667), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(KEYINPUT47), .Z(new_n922));
  OAI21_X1  g497(.A(new_n916), .B1(new_n667), .B2(new_n735), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n667), .B2(new_n737), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n699), .B(new_n702), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(new_n915), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n579), .A2(new_n706), .A3(new_n914), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT48), .Z(new_n929));
  NOR2_X1   g504(.A1(new_n752), .A2(G2067), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n697), .A2(new_n698), .A3(new_n702), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n927), .A2(new_n929), .B1(new_n915), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n922), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(G305), .A2(G1981), .ZN(new_n935));
  INV_X1    g510(.A(G86), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n571), .B1(new_n936), .B2(new_n554), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G1981), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G8), .ZN(new_n942));
  INV_X1    g517(.A(new_n913), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n494), .A2(new_n496), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n488), .A2(new_n491), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n935), .B(new_n938), .C1(KEYINPUT116), .C2(KEYINPUT49), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1976), .ZN(new_n950));
  INV_X1    g525(.A(G288), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n935), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT115), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n913), .B1(new_n946), .B2(new_n954), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n957), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n792), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n913), .B1(new_n965), .B2(new_n912), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n964), .B(new_n911), .C1(G164), .C2(G1384), .ZN(new_n967));
  AOI21_X1  g542(.A(G1971), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G303), .A2(G8), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n972));
  OAI221_X1 g547(.A(G8), .B1(new_n962), .B2(new_n968), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n951), .A2(G1976), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n947), .B1(G288), .B2(new_n950), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT52), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(KEYINPUT52), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n949), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n953), .A2(new_n947), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n973), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n971), .A2(new_n972), .ZN(new_n982));
  OAI21_X1  g557(.A(G8), .B1(new_n962), .B2(new_n968), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n963), .A2(new_n912), .A3(new_n943), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n959), .A2(G2084), .B1(new_n985), .B2(G1966), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT63), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n987), .A2(new_n988), .A3(G286), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n981), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n944), .A2(new_n945), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n954), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n994), .A3(new_n943), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n968), .B1(new_n792), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n982), .B1(new_n997), .B2(new_n942), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n987), .A2(G286), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n979), .A2(new_n998), .A3(new_n973), .A4(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n1000), .A2(new_n988), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n980), .B1(new_n990), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(G2078), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1003), .A2(new_n959), .B1(new_n985), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n911), .B(G1384), .C1(new_n944), .C2(new_n945), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n912), .B1(new_n1007), .B2(KEYINPUT114), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1008), .A2(new_n780), .A3(new_n967), .A4(new_n943), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1009), .A2(KEYINPUT123), .A3(new_n1004), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT123), .B1(new_n1009), .B2(new_n1004), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G171), .ZN(new_n1013));
  OAI211_X1 g588(.A(G301), .B(new_n1006), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(KEYINPUT54), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT126), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1013), .A2(KEYINPUT126), .A3(KEYINPUT54), .A4(new_n1014), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1008), .A2(new_n967), .A3(new_n943), .A4(new_n1020), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT117), .B(G1956), .C1(new_n956), .C2(new_n991), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n995), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n557), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n561), .A2(G91), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(new_n551), .A3(KEYINPUT57), .A4(new_n553), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n959), .A2(new_n743), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n943), .A2(new_n946), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(G2067), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n593), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n1021), .C1(new_n1022), .C2(new_n1025), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(KEYINPUT118), .A3(new_n1039), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1035), .A2(KEYINPUT60), .A3(new_n592), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1032), .A2(new_n592), .A3(new_n1034), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1036), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(KEYINPUT60), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n995), .A2(new_n1024), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT117), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n995), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1038), .B1(new_n1052), .B2(new_n1021), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1039), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1031), .A2(KEYINPUT61), .A3(new_n1039), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1047), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1008), .A2(new_n667), .A3(new_n967), .A4(new_n943), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  AOI22_X1  g636(.A1(new_n1059), .A2(new_n1060), .B1(new_n1033), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n966), .A2(KEYINPUT119), .A3(new_n667), .A4(new_n967), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n543), .A2(KEYINPUT120), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1058), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g642(.A(KEYINPUT59), .B(new_n1065), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1042), .B(new_n1043), .C1(new_n1057), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n985), .A2(new_n1005), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n960), .B2(G1961), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1009), .A2(new_n1004), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1009), .A2(KEYINPUT123), .A3(new_n1004), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1071), .B1(new_n1078), .B2(G301), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1012), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1014), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(KEYINPUT125), .A3(G301), .A4(new_n1006), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n987), .B(KEYINPUT51), .C1(new_n942), .C2(G168), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n986), .A2(G8), .A3(new_n881), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(G8), .C1(new_n986), .C2(new_n881), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT121), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1094), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1019), .A2(new_n1070), .A3(new_n1087), .A4(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1093), .A2(new_n1100), .A3(new_n1095), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n981), .A2(new_n998), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1002), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n579), .B(G1986), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n915), .B1(new_n926), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n934), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT127), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT127), .B(new_n934), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g687(.A1(G319), .A2(new_n636), .ZN(new_n1114));
  NOR3_X1   g688(.A1(G229), .A2(G227), .A3(new_n1114), .ZN(new_n1115));
  OAI211_X1 g689(.A(new_n839), .B(new_n1115), .C1(new_n907), .C2(new_n908), .ZN(G225));
  INV_X1    g690(.A(G225), .ZN(G308));
endmodule


