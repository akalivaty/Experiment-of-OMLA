

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U555 ( .A1(G160), .A2(G40), .ZN(n768) );
  NAND2_X2 U556 ( .A1(n690), .A2(n769), .ZN(n733) );
  AND2_X1 U557 ( .A1(n707), .A2(n700), .ZN(n701) );
  INV_X1 U558 ( .A(G2105), .ZN(n555) );
  AND2_X1 U559 ( .A1(n978), .A2(n812), .ZN(n523) );
  NOR2_X2 U560 ( .A1(n568), .A2(n567), .ZN(G160) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n717) );
  XNOR2_X1 U562 ( .A(n718), .B(n717), .ZN(n723) );
  NOR2_X1 U563 ( .A1(n798), .A2(n523), .ZN(n799) );
  NOR2_X1 U564 ( .A1(n641), .A2(G651), .ZN(n651) );
  XNOR2_X1 U565 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n530) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n524) );
  XNOR2_X1 U567 ( .A(n524), .B(KEYINPUT64), .ZN(n656) );
  NAND2_X1 U568 ( .A1(G89), .A2(n656), .ZN(n525) );
  XNOR2_X1 U569 ( .A(n525), .B(KEYINPUT4), .ZN(n527) );
  XOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  INV_X1 U571 ( .A(G651), .ZN(n531) );
  NOR2_X1 U572 ( .A1(n641), .A2(n531), .ZN(n655) );
  NAND2_X1 U573 ( .A1(G76), .A2(n655), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n528), .B(KEYINPUT5), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n530), .B(n529), .ZN(n539) );
  NOR2_X1 U577 ( .A1(G543), .A2(n531), .ZN(n533) );
  XNOR2_X1 U578 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n532) );
  XNOR2_X1 U579 ( .A(n533), .B(n532), .ZN(n650) );
  NAND2_X1 U580 ( .A1(G63), .A2(n650), .ZN(n535) );
  NAND2_X1 U581 ( .A1(G51), .A2(n651), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U583 ( .A(n536), .B(KEYINPUT6), .ZN(n537) );
  XNOR2_X1 U584 ( .A(KEYINPUT78), .B(n537), .ZN(n538) );
  NOR2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U586 ( .A(KEYINPUT7), .B(n540), .Z(G168) );
  XNOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .ZN(n541) );
  XNOR2_X1 U588 ( .A(n541), .B(KEYINPUT79), .ZN(G286) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G57), .ZN(G237) );
  INV_X1 U591 ( .A(G69), .ZN(G235) );
  INV_X1 U592 ( .A(G108), .ZN(G238) );
  INV_X1 U593 ( .A(G120), .ZN(G236) );
  INV_X1 U594 ( .A(G132), .ZN(G219) );
  INV_X1 U595 ( .A(G82), .ZN(G220) );
  NAND2_X1 U596 ( .A1(G52), .A2(n651), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT69), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n655), .A2(G77), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G90), .A2(n656), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U601 ( .A(n545), .B(KEYINPUT9), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G64), .A2(n650), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U605 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U606 ( .A1(n887), .A2(G114), .ZN(n550) );
  XOR2_X1 U607 ( .A(KEYINPUT91), .B(n550), .Z(n552) );
  NOR2_X1 U608 ( .A1(G2104), .A2(n555), .ZN(n884) );
  NAND2_X1 U609 ( .A1(n884), .A2(G126), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT92), .ZN(n560) );
  NOR2_X1 U612 ( .A1(G2104), .A2(G2105), .ZN(n554) );
  XOR2_X1 U613 ( .A(KEYINPUT17), .B(n554), .Z(n879) );
  NAND2_X1 U614 ( .A1(G138), .A2(n879), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n555), .A2(G2104), .ZN(n556) );
  XNOR2_X2 U616 ( .A(n556), .B(KEYINPUT65), .ZN(n880) );
  NAND2_X1 U617 ( .A1(G102), .A2(n880), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U619 ( .A1(n560), .A2(n559), .ZN(G164) );
  NAND2_X1 U620 ( .A1(G125), .A2(n884), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G137), .A2(n879), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G113), .A2(n887), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT66), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G101), .A2(n880), .ZN(n564) );
  XOR2_X1 U626 ( .A(n564), .B(KEYINPUT23), .Z(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U629 ( .A(n569), .B(KEYINPUT10), .Z(n917) );
  NAND2_X1 U630 ( .A1(n917), .A2(G567), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n650), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U634 ( .A1(G81), .A2(n656), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G68), .A2(n655), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n651), .A2(G43), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n982) );
  INV_X1 U642 ( .A(G860), .ZN(n603) );
  NOR2_X1 U643 ( .A1(n982), .A2(n603), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT72), .B(n580), .Z(G153) );
  INV_X1 U645 ( .A(G171), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U647 ( .A1(G66), .A2(n650), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G92), .A2(n656), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT73), .B(n583), .Z(n589) );
  NAND2_X1 U651 ( .A1(n655), .A2(G79), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(KEYINPUT74), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G54), .A2(n651), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U655 ( .A(KEYINPUT75), .B(n587), .Z(n588) );
  NOR2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U657 ( .A(KEYINPUT15), .B(n590), .ZN(n708) );
  INV_X1 U658 ( .A(G868), .ZN(n672) );
  NAND2_X1 U659 ( .A1(n708), .A2(n672), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U661 ( .A1(n650), .A2(G65), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n655), .A2(G78), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G91), .A2(n656), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n651), .A2(G53), .ZN(n595) );
  XOR2_X1 U666 ( .A(KEYINPUT70), .B(n595), .Z(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U669 ( .A(KEYINPUT71), .B(n600), .ZN(n972) );
  INV_X1 U670 ( .A(n972), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G286), .A2(G868), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G299), .A2(n672), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U675 ( .A(n708), .ZN(n987) );
  NAND2_X1 U676 ( .A1(n604), .A2(n987), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n982), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G868), .A2(n987), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n884), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n887), .A2(G111), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G135), .A2(n879), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G99), .A2(n880), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n919) );
  XOR2_X1 U690 ( .A(G2096), .B(n919), .Z(n616) );
  NOR2_X1 U691 ( .A1(G2100), .A2(n616), .ZN(n617) );
  XOR2_X1 U692 ( .A(KEYINPUT80), .B(n617), .Z(G156) );
  NAND2_X1 U693 ( .A1(G67), .A2(n650), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G93), .A2(n656), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G80), .A2(n655), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT81), .B(n620), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n651), .A2(G55), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n671) );
  NAND2_X1 U701 ( .A1(G559), .A2(n987), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(n982), .ZN(n669) );
  NOR2_X1 U703 ( .A1(G860), .A2(n669), .ZN(n626) );
  XOR2_X1 U704 ( .A(n671), .B(n626), .Z(G145) );
  NAND2_X1 U705 ( .A1(G85), .A2(n656), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n650), .A2(G60), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G72), .A2(n655), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G47), .A2(n651), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT68), .B(n633), .Z(G290) );
  NAND2_X1 U713 ( .A1(G61), .A2(n650), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G86), .A2(n656), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n655), .A2(G73), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n651), .A2(G48), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G87), .A2(n641), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G651), .A2(G74), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(KEYINPUT82), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G49), .A2(n651), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U726 ( .A1(n650), .A2(n645), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT83), .B(n646), .Z(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT84), .ZN(G288) );
  NAND2_X1 U730 ( .A1(G62), .A2(n650), .ZN(n653) );
  NAND2_X1 U731 ( .A1(G50), .A2(n651), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(KEYINPUT85), .B(n654), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n655), .A2(G75), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G88), .A2(n656), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U737 ( .A(KEYINPUT86), .B(n659), .Z(n660) );
  NAND2_X1 U738 ( .A1(n661), .A2(n660), .ZN(G303) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n663) );
  XNOR2_X1 U741 ( .A(G305), .B(KEYINPUT88), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U743 ( .A(n664), .B(G288), .Z(n666) );
  XOR2_X1 U744 ( .A(G299), .B(G166), .Z(n665) );
  XNOR2_X1 U745 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U746 ( .A(G290), .B(n667), .Z(n668) );
  XNOR2_X1 U747 ( .A(n671), .B(n668), .ZN(n897) );
  XNOR2_X1 U748 ( .A(n669), .B(n897), .ZN(n670) );
  NAND2_X1 U749 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U750 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U752 ( .A(KEYINPUT89), .B(n675), .Z(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U761 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G96), .A2(n682), .ZN(n821) );
  NAND2_X1 U763 ( .A1(n821), .A2(G2106), .ZN(n687) );
  NOR2_X1 U764 ( .A1(G236), .A2(G238), .ZN(n684) );
  NOR2_X1 U765 ( .A1(G235), .A2(G237), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U767 ( .A(KEYINPUT90), .B(n685), .ZN(n822) );
  NAND2_X1 U768 ( .A1(n822), .A2(G567), .ZN(n686) );
  NAND2_X1 U769 ( .A1(n687), .A2(n686), .ZN(n823) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n823), .A2(n688), .ZN(n820) );
  NAND2_X1 U772 ( .A1(n820), .A2(G36), .ZN(G176) );
  INV_X1 U773 ( .A(KEYINPUT96), .ZN(n689) );
  XNOR2_X1 U774 ( .A(n768), .B(n689), .ZN(n690) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U776 ( .A1(G8), .A2(n733), .ZN(n761) );
  NOR2_X1 U777 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U778 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  NOR2_X1 U779 ( .A1(n761), .A2(n692), .ZN(n766) );
  INV_X1 U780 ( .A(n733), .ZN(n719) );
  NAND2_X1 U781 ( .A1(n719), .A2(G2072), .ZN(n693) );
  XNOR2_X1 U782 ( .A(n693), .B(KEYINPUT27), .ZN(n695) );
  INV_X1 U783 ( .A(G1956), .ZN(n837) );
  NOR2_X1 U784 ( .A1(n837), .A2(n719), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n712) );
  NOR2_X1 U786 ( .A1(n972), .A2(n712), .ZN(n696) );
  XOR2_X1 U787 ( .A(n696), .B(KEYINPUT28), .Z(n716) );
  INV_X1 U788 ( .A(n733), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n697), .A2(G1996), .ZN(n698) );
  XOR2_X1 U790 ( .A(KEYINPUT26), .B(n698), .Z(n699) );
  NOR2_X2 U791 ( .A1(n982), .A2(n699), .ZN(n707) );
  NAND2_X1 U792 ( .A1(G1341), .A2(n733), .ZN(n706) );
  AND2_X1 U793 ( .A1(n706), .A2(n987), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n701), .B(KEYINPUT97), .ZN(n705) );
  NOR2_X1 U795 ( .A1(n719), .A2(G1348), .ZN(n703) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n733), .ZN(n702) );
  NOR2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n972), .A2(n712), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n718) );
  OR2_X1 U805 ( .A1(n719), .A2(G1961), .ZN(n721) );
  XNOR2_X1 U806 ( .A(KEYINPUT25), .B(G2078), .ZN(n951) );
  NAND2_X1 U807 ( .A1(n719), .A2(n951), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n727), .A2(G171), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n732) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n761), .ZN(n744) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n733), .ZN(n741) );
  NOR2_X1 U813 ( .A1(n744), .A2(n741), .ZN(n724) );
  NAND2_X1 U814 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U816 ( .A1(G168), .A2(n726), .ZN(n729) );
  NOR2_X1 U817 ( .A1(G171), .A2(n727), .ZN(n728) );
  NOR2_X1 U818 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(n730), .Z(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n742) );
  NAND2_X1 U821 ( .A1(n742), .A2(G286), .ZN(n738) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n761), .ZN(n735) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G8), .A2(n739), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n740), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U829 ( .A1(G8), .A2(n741), .ZN(n746) );
  INV_X1 U830 ( .A(n742), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n760) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n753), .A2(n749), .ZN(n976) );
  NAND2_X1 U837 ( .A1(n760), .A2(n976), .ZN(n750) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NAND2_X1 U839 ( .A1(n750), .A2(n980), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n761), .A2(n751), .ZN(n752) );
  NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n752), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n754), .A2(n761), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n969) );
  NAND2_X1 U846 ( .A1(n757), .A2(n969), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  INV_X1 U853 ( .A(n767), .ZN(n800) );
  NOR2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n812) );
  XOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .Z(n770) );
  XNOR2_X1 U856 ( .A(KEYINPUT93), .B(n770), .ZN(n801) );
  NAND2_X1 U857 ( .A1(n880), .A2(G104), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n771), .B(KEYINPUT94), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G140), .A2(n879), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G116), .A2(n887), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G128), .A2(n884), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n780), .ZN(n856) );
  NOR2_X1 U868 ( .A1(n801), .A2(n856), .ZN(n933) );
  NAND2_X1 U869 ( .A1(n812), .A2(n933), .ZN(n809) );
  NAND2_X1 U870 ( .A1(G131), .A2(n879), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G95), .A2(n880), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G107), .A2(n887), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G119), .A2(n884), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n866) );
  INV_X1 U877 ( .A(G1991), .ZN(n832) );
  NOR2_X1 U878 ( .A1(n866), .A2(n832), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G105), .A2(n880), .ZN(n787) );
  XNOR2_X1 U880 ( .A(n787), .B(KEYINPUT38), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G117), .A2(n887), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G129), .A2(n884), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G141), .A2(n879), .ZN(n790) );
  XNOR2_X1 U885 ( .A(KEYINPUT95), .B(n790), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n855) );
  AND2_X1 U888 ( .A1(n855), .A2(G1996), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n931) );
  INV_X1 U890 ( .A(n931), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n797), .A2(n812), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n809), .A2(n802), .ZN(n798) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n815) );
  NAND2_X1 U895 ( .A1(n801), .A2(n856), .ZN(n942) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n855), .ZN(n926) );
  INV_X1 U897 ( .A(n802), .ZN(n806) );
  AND2_X1 U898 ( .A1(n832), .A2(n866), .ZN(n803) );
  XNOR2_X1 U899 ( .A(KEYINPUT98), .B(n803), .ZN(n918) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n918), .A2(n804), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n926), .A2(n807), .ZN(n808) );
  XNOR2_X1 U904 ( .A(KEYINPUT39), .B(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n942), .A2(n811), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n917), .ZN(G217) );
  NAND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT100), .B(n817), .Z(n818) );
  NAND2_X1 U913 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(G188) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  INV_X1 U920 ( .A(n823), .ZN(G319) );
  XOR2_X1 U921 ( .A(G2100), .B(G2096), .Z(n825) );
  XNOR2_X1 U922 ( .A(KEYINPUT42), .B(G2678), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(G2090), .Z(n827) );
  XNOR2_X1 U925 ( .A(G2067), .B(G2072), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U927 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U928 ( .A(G2078), .B(G2084), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(G227) );
  XOR2_X1 U930 ( .A(G1976), .B(G1971), .Z(n834) );
  XOR2_X1 U931 ( .A(G1996), .B(n832), .Z(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n845) );
  XOR2_X1 U933 ( .A(KEYINPUT103), .B(G2474), .Z(n836) );
  XNOR2_X1 U934 ( .A(G1981), .B(KEYINPUT101), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n837), .B(G1961), .ZN(n839) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT41), .B(KEYINPUT102), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(n845), .B(n844), .Z(G229) );
  NAND2_X1 U943 ( .A1(G124), .A2(n884), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n846), .B(KEYINPUT104), .ZN(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT44), .B(n847), .ZN(n850) );
  NAND2_X1 U946 ( .A1(G112), .A2(n887), .ZN(n848) );
  XOR2_X1 U947 ( .A(KEYINPUT105), .B(n848), .Z(n849) );
  NAND2_X1 U948 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U949 ( .A1(G136), .A2(n879), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G100), .A2(n880), .ZN(n851) );
  NAND2_X1 U951 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U952 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U953 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U954 ( .A(G164), .B(G160), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n865) );
  XOR2_X1 U956 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n860) );
  XNOR2_X1 U957 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n861), .B(KEYINPUT46), .Z(n863) );
  XNOR2_X1 U960 ( .A(n919), .B(KEYINPUT107), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U962 ( .A(n865), .B(n864), .Z(n868) );
  XNOR2_X1 U963 ( .A(n866), .B(G162), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n868), .B(n867), .ZN(n893) );
  NAND2_X1 U965 ( .A1(n880), .A2(G103), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n869), .B(KEYINPUT108), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G139), .A2(n879), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n878) );
  NAND2_X1 U969 ( .A1(n884), .A2(G127), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT109), .B(n872), .Z(n874) );
  NAND2_X1 U971 ( .A1(n887), .A2(G115), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT110), .B(n876), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n935) );
  NAND2_X1 U976 ( .A1(G142), .A2(n879), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G106), .A2(n880), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n883), .B(KEYINPUT45), .ZN(n886) );
  NAND2_X1 U980 ( .A1(G130), .A2(n884), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n890) );
  NAND2_X1 U982 ( .A1(n887), .A2(G118), .ZN(n888) );
  XOR2_X1 U983 ( .A(KEYINPUT106), .B(n888), .Z(n889) );
  NOR2_X1 U984 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U985 ( .A(n935), .B(n891), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U987 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n982), .B(KEYINPUT114), .ZN(n896) );
  XOR2_X1 U989 ( .A(G301), .B(n987), .Z(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n899) );
  XOR2_X1 U991 ( .A(n897), .B(G286), .Z(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U993 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U994 ( .A(G2454), .B(G2435), .Z(n902) );
  XNOR2_X1 U995 ( .A(G2438), .B(G2427), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n909) );
  XOR2_X1 U997 ( .A(KEYINPUT99), .B(G2446), .Z(n904) );
  XNOR2_X1 U998 ( .A(G2443), .B(G2430), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n905), .B(G2451), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(n910), .A2(G14), .ZN(n916) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n916), .ZN(G401) );
  INV_X1 U1013 ( .A(n917), .ZN(G223) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1015 ( .A(KEYINPUT115), .B(n920), .Z(n922) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(KEYINPUT116), .B(n923), .ZN(n929) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G162), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(KEYINPUT117), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT51), .B(n927), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1026 ( .A(KEYINPUT118), .B(n934), .Z(n940) );
  XOR2_X1 U1027 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1032 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1033 ( .A(n943), .B(KEYINPUT52), .ZN(n944) );
  XNOR2_X1 U1034 ( .A(KEYINPUT119), .B(n944), .ZN(n946) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1037 ( .A1(n947), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1038 ( .A(G2090), .B(G35), .ZN(n960) );
  XOR2_X1 U1039 ( .A(G25), .B(G1991), .Z(n948) );
  NAND2_X1 U1040 ( .A1(n948), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n955) );
  XOR2_X1 U1044 ( .A(n951), .B(G27), .Z(n953) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1054 ( .A(KEYINPUT55), .B(n964), .Z(n966) );
  INV_X1 U1055 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n967), .ZN(n1025) );
  XOR2_X1 U1058 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n968) );
  XOR2_X1 U1059 ( .A(G16), .B(n968), .Z(n993) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(KEYINPUT57), .ZN(n991) );
  XOR2_X1 U1063 ( .A(n972), .B(G1956), .Z(n974) );
  AND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(n981), .B(KEYINPUT121), .ZN(n986) );
  XOR2_X1 U1070 ( .A(G171), .B(G1961), .Z(n984) );
  XNOR2_X1 U1071 ( .A(n982), .B(G1341), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1074 ( .A(G1348), .B(n987), .Z(n988) );
  NOR2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1077 ( .A1(n993), .A2(n992), .ZN(n1023) );
  INV_X1 U1078 ( .A(G16), .ZN(n1021) );
  XOR2_X1 U1079 ( .A(G5), .B(G1961), .Z(n1016) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1976), .B(G23), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(KEYINPUT126), .B(n996), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1986), .B(KEYINPUT127), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n997), .B(G24), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(n1000), .B(KEYINPUT58), .ZN(n1014) );
  XOR2_X1 U1088 ( .A(G20), .B(G1956), .Z(n1003) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT122), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1006), .Z(n1010) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT124), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G1348), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT60), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT125), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(G21), .B(G1966), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .ZN(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

