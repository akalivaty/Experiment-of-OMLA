//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  XOR2_X1   g045(.A(new_n470), .B(KEYINPUT71), .Z(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n469), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n475), .A2(new_n476), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n473), .A2(new_n469), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(KEYINPUT73), .B2(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n468), .A2(new_n469), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n477), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n468), .A2(KEYINPUT72), .A3(G126), .A4(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n473), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n496), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT74), .B1(new_n509), .B2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(new_n507), .A3(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(KEYINPUT75), .A3(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n506), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n507), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n524), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n510), .A2(new_n512), .ZN(new_n529));
  INV_X1    g104(.A(new_n508), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n529), .A2(G51), .A3(G543), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n514), .A2(KEYINPUT75), .A3(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT75), .B1(new_n514), .B2(G543), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT76), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n513), .A2(new_n520), .A3(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n531), .A2(KEYINPUT76), .A3(new_n536), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n538), .A2(new_n542), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(new_n520), .A2(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n507), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n513), .A2(new_n520), .A3(G90), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n513), .A2(G52), .A3(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT77), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n548), .B1(new_n552), .B2(new_n554), .ZN(G171));
  AOI22_X1  g130(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n507), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n513), .A2(new_n520), .A3(G81), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n513), .A2(G43), .A3(G543), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n560), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n520), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n521), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G91), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n530), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(KEYINPUT79), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n513), .A2(new_n585), .A3(G53), .A4(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(KEYINPUT9), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n578), .A2(new_n580), .A3(new_n583), .A4(new_n587), .ZN(G299));
  AND3_X1   g163(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n553), .B1(new_n549), .B2(new_n550), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n546), .A2(new_n547), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n589), .A2(new_n590), .B1(new_n507), .B2(new_n591), .ZN(G301));
  OAI21_X1  g167(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT81), .ZN(new_n594));
  INV_X1    g169(.A(new_n522), .ZN(new_n595));
  AOI22_X1  g170(.A1(G87), .A2(new_n579), .B1(new_n595), .B2(G49), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT82), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G288));
  AND3_X1   g174(.A1(new_n513), .A2(new_n520), .A3(G86), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT83), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n507), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(G48), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(KEYINPUT83), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n601), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(G305));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  INV_X1    g182(.A(G47), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n607), .A2(new_n521), .B1(new_n522), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n507), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n609), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n595), .A2(G54), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n513), .A2(new_n520), .A3(G92), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n513), .A2(new_n520), .A3(new_n617), .A4(G92), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n572), .B2(new_n574), .ZN(new_n623));
  AND2_X1   g198(.A1(G79), .A2(G543), .ZN(new_n624));
  OAI21_X1  g199(.A(G651), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n626));
  AND4_X1   g201(.A1(new_n614), .A2(new_n621), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n613), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n613), .B1(new_n627), .B2(G868), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n468), .A2(new_n478), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n483), .A2(G135), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT86), .ZN(new_n646));
  INV_X1    g221(.A(G111), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n476), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n482), .A2(G123), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(G2096), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n642), .A2(new_n643), .ZN(new_n657));
  INV_X1    g232(.A(new_n654), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G2096), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n644), .A2(new_n656), .A3(new_n657), .A4(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT88), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2427), .B(G2430), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(KEYINPUT14), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(G401));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n643), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n680), .B2(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n655), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n693), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n697), .B(new_n698), .S(new_n691), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1971), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n707), .A2(G23), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n597), .B2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT33), .B(G1976), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n707), .A2(G6), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G305), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(new_n714), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n715), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n717), .A2(new_n719), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n710), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n707), .A2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G290), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n707), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT90), .Z(new_n735));
  AOI22_X1  g310(.A1(G119), .A2(new_n482), .B1(new_n483), .B2(G131), .ZN(new_n736));
  OAI221_X1 g311(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n726), .A2(new_n727), .A3(new_n732), .A4(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(KEYINPUT36), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(KEYINPUT92), .ZN(new_n747));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n743), .B2(KEYINPUT36), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n745), .A2(KEYINPUT36), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n744), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n733), .A2(G32), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n482), .A2(G129), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n751), .B1(new_n761), .B2(new_n733), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT27), .ZN(new_n763));
  INV_X1    g338(.A(G1996), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n733), .A2(G33), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n483), .A2(G139), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n770), .C1(new_n469), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(KEYINPUT24), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(KEYINPUT24), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(KEYINPUT95), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(KEYINPUT95), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n480), .B2(new_n733), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n766), .A2(new_n773), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n733), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n783), .B(new_n784), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n482), .A2(G128), .ZN(new_n786));
  OAI221_X1 g361(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n483), .A2(G140), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n785), .B1(new_n789), .B2(new_n733), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n781), .B(new_n791), .C1(new_n766), .C2(new_n773), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n733), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n733), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT29), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G2090), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT31), .B(G11), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(G28), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n733), .B1(new_n799), .B2(G28), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n798), .B1(new_n800), .B2(new_n801), .C1(new_n658), .C2(new_n733), .ZN(new_n802));
  INV_X1    g377(.A(G2078), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n504), .A2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n733), .A2(G27), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n802), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n806), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n808), .A2(G2078), .B1(new_n780), .B2(new_n779), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n792), .A2(new_n796), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n765), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n707), .A2(G19), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n564), .B2(new_n707), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1341), .Z(new_n814));
  INV_X1    g389(.A(G1348), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n627), .A2(new_n707), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G4), .B2(new_n707), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g394(.A1(G168), .A2(new_n707), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n707), .B2(G21), .ZN(new_n821));
  INV_X1    g396(.A(G1966), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT98), .ZN(new_n824));
  NOR2_X1   g399(.A1(G171), .A2(new_n707), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G5), .B2(new_n707), .ZN(new_n826));
  INV_X1    g401(.A(G1961), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n821), .A2(new_n822), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n811), .A2(new_n819), .A3(new_n824), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n795), .A2(G2090), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT99), .Z(new_n832));
  XOR2_X1   g407(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n707), .A2(G20), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n631), .B2(new_n707), .ZN(new_n836));
  INV_X1    g411(.A(G1956), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT101), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n747), .A2(new_n750), .A3(new_n842), .ZN(G311));
  INV_X1    g418(.A(new_n747), .ZN(new_n844));
  INV_X1    g419(.A(new_n750), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n841), .ZN(G150));
  NAND2_X1  g421(.A1(new_n520), .A2(G67), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n507), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n595), .A2(G55), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n579), .A2(G93), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(KEYINPUT102), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n855), .A2(new_n521), .B1(new_n522), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n854), .B1(new_n857), .B2(new_n849), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n563), .A2(new_n853), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n558), .A2(new_n559), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT78), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n857), .A2(new_n849), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT102), .A4(new_n557), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT38), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n627), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  INV_X1    g445(.A(G860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n864), .A2(new_n871), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(G145));
  INV_X1    g451(.A(new_n789), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n760), .B(new_n877), .ZN(new_n878));
  OAI221_X1 g453(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n482), .A2(G130), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n483), .A2(new_n881), .A3(G142), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n483), .B2(G142), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n879), .B(new_n880), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n878), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n772), .B(new_n504), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n738), .B(new_n641), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n885), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n480), .B(G162), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n654), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g470(.A(new_n636), .B(new_n866), .Z(new_n896));
  XOR2_X1   g471(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n587), .A2(new_n583), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(KEYINPUT104), .A3(new_n578), .A4(new_n580), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n627), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n621), .A2(new_n625), .A3(new_n614), .A4(new_n626), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(G299), .A3(new_n898), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n897), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n902), .A2(new_n906), .A3(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n896), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n904), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n909), .B2(new_n896), .ZN(new_n910));
  XNOR2_X1  g485(.A(G305), .B(new_n597), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(G290), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n914), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g496(.A(new_n920), .B1(G868), .B2(new_n864), .ZN(G331));
  NAND3_X1  g497(.A1(new_n543), .A2(new_n541), .A3(new_n539), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT107), .B1(new_n923), .B2(new_n537), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n538), .A2(new_n542), .A3(new_n925), .A4(new_n543), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(G171), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(G301), .A2(G286), .A3(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(new_n866), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n907), .B2(new_n905), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n929), .A2(new_n866), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n927), .A2(new_n928), .B1(new_n859), .B2(new_n865), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n904), .A3(new_n902), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n913), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT41), .B1(new_n902), .B2(new_n904), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n940), .B(new_n930), .C1(new_n909), .C2(new_n897), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n913), .B1(new_n941), .B2(new_n935), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT109), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n897), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n902), .A2(new_n904), .A3(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n945), .A2(new_n934), .A3(new_n939), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n930), .A2(new_n909), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n914), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n937), .A4(new_n936), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(KEYINPUT43), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n913), .B1(new_n931), .B2(new_n935), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n938), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(KEYINPUT44), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n938), .B2(new_n952), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n948), .A2(new_n957), .A3(new_n937), .A4(new_n936), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI211_X1 g536(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n956), .C2(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n954), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT110), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(new_n954), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n504), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n471), .A2(G40), .A3(new_n479), .ZN(new_n972));
  OR3_X1    g547(.A1(new_n971), .A2(KEYINPUT111), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT111), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n789), .B(G2067), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n761), .B2(new_n764), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n738), .B(new_n741), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n973), .A2(new_n764), .A3(new_n974), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n973), .A2(new_n985), .A3(new_n764), .A4(new_n974), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n761), .ZN(new_n988));
  XNOR2_X1  g563(.A(G290), .B(G1986), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n973), .A2(new_n974), .A3(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n980), .A2(new_n982), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT114), .Z(new_n992));
  XOR2_X1   g567(.A(KEYINPUT116), .B(G8), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n498), .A2(new_n503), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n995), .B2(new_n496), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n471), .A2(G40), .A3(new_n479), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n996), .B2(new_n997), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n999), .A2(new_n1001), .A3(G2084), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n972), .B1(new_n969), .B2(new_n970), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(KEYINPUT45), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1966), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n994), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G286), .A2(new_n994), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1000), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n969), .A2(new_n970), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n822), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n972), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(new_n780), .A3(new_n998), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1018), .B2(new_n1009), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n993), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1010), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT122), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1011), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1009), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1000), .A2(new_n996), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n994), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n597), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT117), .B(G1976), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n598), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1029), .A3(new_n1037), .A4(new_n994), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1033), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n603), .A2(new_n604), .ZN(new_n1041));
  OAI21_X1  g616(.A(G1981), .B1(new_n1041), .B2(new_n600), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT49), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n1030), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT115), .B(G2090), .Z(new_n1047));
  AND3_X1   g622(.A1(new_n1016), .A2(new_n998), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n994), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1052), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1054), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1046), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n971), .A2(new_n1004), .A3(new_n803), .A4(new_n1000), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n827), .B1(new_n999), .B2(new_n1001), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1003), .A2(KEYINPUT53), .A3(new_n803), .A4(new_n1004), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1062), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT123), .B1(new_n1062), .B2(G171), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1056), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1026), .A2(new_n1028), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT124), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1026), .A2(new_n1068), .A3(new_n1028), .A4(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g645(.A(G286), .B(new_n993), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1046), .A2(new_n1053), .A3(new_n1055), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT118), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1006), .A2(new_n1073), .A3(G286), .ZN(new_n1078));
  OAI21_X1  g653(.A(G8), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1052), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1055), .A3(new_n1046), .A4(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1031), .B(new_n598), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1030), .B1(new_n1083), .B2(new_n1040), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1055), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1046), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT119), .B(G1996), .Z(new_n1088));
  INV_X1    g663(.A(new_n1029), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1087), .A2(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n564), .A2(KEYINPUT120), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(KEYINPUT59), .A3(new_n1093), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1348), .B1(new_n1016), .B2(new_n998), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1029), .A2(G2067), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n903), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1103), .A2(new_n627), .A3(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1003), .A2(new_n1004), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1956), .B1(new_n1016), .B2(new_n998), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n631), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1108), .A2(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n837), .B1(new_n999), .B2(new_n1001), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1107), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1114), .B(new_n1115), .C1(new_n1087), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT61), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1102), .A2(new_n1106), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT61), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1113), .B1(new_n903), .B2(new_n1100), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(new_n1122), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1062), .A2(G171), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(new_n1127), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1062), .A2(G171), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT54), .B1(new_n1129), .B2(new_n1125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1056), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1082), .B(new_n1086), .C1(new_n1124), .C2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n992), .B1(new_n1070), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT47), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT46), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n984), .A2(new_n1137), .A3(new_n986), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT125), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n984), .A2(new_n1140), .A3(new_n1137), .A4(new_n986), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n761), .A2(new_n978), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n977), .A2(new_n1144), .B1(new_n987), .B2(KEYINPUT46), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1143), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1136), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n973), .A2(new_n731), .A3(new_n729), .A4(new_n974), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT48), .ZN(new_n1151));
  AND4_X1   g726(.A1(new_n988), .A2(new_n980), .A3(new_n982), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n738), .A2(new_n741), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n980), .A2(new_n988), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(G2067), .B2(new_n877), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n1155), .B2(new_n977), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT126), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(KEYINPUT47), .A3(new_n1146), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1149), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1135), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g736(.A1(G401), .A2(new_n464), .A3(G227), .ZN(new_n1163));
  AOI211_X1 g737(.A(G229), .B(new_n1163), .C1(new_n892), .C2(new_n893), .ZN(new_n1164));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1165));
  AND3_X1   g739(.A1(new_n1164), .A2(new_n1165), .A3(new_n959), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1164), .B2(new_n959), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1167), .ZN(G308));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n959), .ZN(G225));
endmodule


