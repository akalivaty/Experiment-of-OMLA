//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT89), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(KEYINPUT89), .A3(new_n207), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n206), .B2(KEYINPUT88), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n203), .A2(KEYINPUT88), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(KEYINPUT14), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n218), .A2(KEYINPUT14), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(KEYINPUT14), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n222), .B(new_n223), .C1(G29gat), .C2(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n215), .A2(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n226), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n228), .A2(new_n217), .A3(new_n221), .A4(new_n224), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT87), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT17), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  AOI211_X1 g032(.A(KEYINPUT87), .B(new_n233), .C1(new_n227), .C2(new_n229), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n214), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n211), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n212), .A2(new_n213), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n230), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n240), .B(KEYINPUT13), .Z(new_n244));
  INV_X1    g043(.A(new_n239), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n238), .A2(new_n230), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n235), .A2(new_n239), .A3(KEYINPUT18), .A4(new_n240), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT11), .B(G169gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(G113gat), .B(G141gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n243), .A2(new_n247), .A3(new_n254), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT90), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G1gat), .B(G29gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(G127gat), .ZN(new_n269));
  INV_X1    g068(.A(G120gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G113gat), .ZN(new_n271));
  INV_X1    g070(.A(G113gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G120gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI211_X1 g075(.A(KEYINPUT1), .B(G127gat), .C1(new_n271), .C2(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n268), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G162gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G155gat), .ZN(new_n280));
  INV_X1    g079(.A(G155gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(KEYINPUT2), .ZN(new_n285));
  INV_X1    g084(.A(G148gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G155gat), .B(G162gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT2), .B1(new_n292), .B2(new_n281), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  OAI21_X1  g095(.A(G127gat), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n275), .A3(new_n269), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(G134gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n294), .A3(new_n307), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n297), .A2(new_n298), .A3(G134gat), .ZN(new_n309));
  AOI21_X1  g108(.A(G134gat), .B1(new_n297), .B2(new_n298), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n305), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n278), .A2(new_n295), .A3(new_n299), .A4(new_n301), .ZN(new_n312));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n303), .A2(new_n311), .A3(new_n312), .A4(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n317), .B1(new_n300), .B2(new_n313), .ZN(new_n320));
  INV_X1    g119(.A(new_n311), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n300), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT5), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n267), .B(new_n316), .C1(new_n322), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT77), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n300), .A2(new_n313), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n318), .A3(new_n311), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n324), .B2(new_n314), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n303), .A2(new_n311), .A3(new_n312), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n335), .A2(new_n337), .B1(new_n338), .B2(new_n315), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT78), .B1(new_n339), .B2(new_n267), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n316), .B1(new_n322), .B2(new_n326), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342));
  INV_X1    g141(.A(new_n267), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n330), .A2(new_n332), .A3(new_n340), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT79), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n339), .A2(new_n267), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT6), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n340), .A2(new_n344), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n332), .A4(new_n330), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G169gat), .ZN(new_n353));
  INV_X1    g152(.A(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n353), .B2(new_n354), .ZN(new_n357));
  NOR2_X1   g156(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(KEYINPUT24), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n361), .A2(KEYINPUT24), .ZN(new_n363));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT23), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n359), .A2(new_n362), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT25), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT67), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT26), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n355), .A2(KEYINPUT26), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n376), .A3(new_n375), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n374), .A2(new_n379), .A3(new_n381), .A4(new_n361), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n362), .A2(new_n363), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT64), .B(G169gat), .Z(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(KEYINPUT23), .A3(new_n354), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n383), .A2(new_n385), .A3(new_n386), .A4(new_n359), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n367), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT29), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n389), .B2(new_n388), .ZN(new_n393));
  INV_X1    g192(.A(G218gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT70), .ZN(new_n395));
  INV_X1    g194(.A(G211gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(G218gat), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G197gat), .B(G204gat), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n401), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n396), .B1(new_n401), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n394), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT22), .B1(new_n408), .B2(G218gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n402), .ZN(new_n410));
  OAI21_X1  g209(.A(G211gat), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n401), .A2(new_n396), .A3(new_n402), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(G218gat), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n393), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n393), .A2(new_n415), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT71), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G8gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(new_n220), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n416), .B2(new_n417), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n418), .A2(new_n427), .A3(new_n423), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n405), .B2(new_n413), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n304), .B1(new_n432), .B2(new_n306), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n308), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n405), .A2(new_n413), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n403), .A2(new_n404), .A3(new_n394), .ZN(new_n438));
  AOI21_X1  g237(.A(G218gat), .B1(new_n411), .B2(new_n412), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n434), .B(new_n304), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(new_n436), .A3(new_n305), .A4(new_n431), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(G22gat), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n437), .A2(new_n442), .A3(G22gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(KEYINPUT81), .ZN(new_n445));
  XOR2_X1   g244(.A(G78gat), .B(G106gat), .Z(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT31), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n447), .B(G50gat), .Z(new_n448));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n449), .B(G22gat), .C1(new_n437), .C2(new_n442), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n448), .ZN(new_n452));
  INV_X1    g251(.A(G22gat), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n295), .B1(new_n454), .B2(new_n307), .ZN(new_n455));
  INV_X1    g254(.A(new_n436), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n430), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n453), .B1(new_n457), .B2(new_n441), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n452), .B1(new_n444), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(KEYINPUT80), .B(new_n452), .C1(new_n444), .C2(new_n458), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n451), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n278), .A2(new_n299), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n388), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n309), .A2(new_n310), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n467), .A2(new_n367), .A3(new_n387), .A4(new_n382), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT32), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G71gat), .ZN(new_n472));
  INV_X1    g271(.A(G99gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n475));
  AND2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n469), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n470), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n474), .B1(new_n469), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n474), .C1(new_n469), .C2(new_n479), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n468), .A3(new_n464), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT34), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n466), .A2(new_n468), .A3(new_n487), .A4(new_n464), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n489), .B(new_n477), .C1(new_n481), .C2(new_n483), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n352), .A2(new_n429), .A3(new_n463), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n481), .A2(new_n483), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n489), .B1(new_n496), .B2(new_n477), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n484), .A2(new_n490), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(KEYINPUT84), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n491), .B2(new_n492), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n463), .A2(new_n429), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n348), .B(KEYINPUT83), .ZN(new_n503));
  INV_X1    g302(.A(new_n347), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n328), .A4(new_n327), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT82), .B1(new_n329), .B2(new_n347), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT85), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n499), .A2(new_n501), .A3(new_n429), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT35), .B1(new_n503), .B2(new_n508), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n463), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n463), .ZN(new_n518));
  INV_X1    g317(.A(new_n352), .ZN(new_n519));
  INV_X1    g318(.A(new_n429), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR3_X1    g320(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT37), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT37), .B1(new_n416), .B2(new_n417), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n422), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(KEYINPUT38), .ZN(new_n525));
  INV_X1    g324(.A(new_n424), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(KEYINPUT38), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n503), .A2(new_n525), .A3(new_n527), .A4(new_n508), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n338), .A2(new_n313), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(KEYINPUT39), .C1(new_n314), .C2(new_n324), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n267), .C1(KEYINPUT39), .C2(new_n529), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT40), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n520), .A2(new_n504), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n528), .B(new_n463), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n493), .B(KEYINPUT36), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n260), .B1(new_n517), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G71gat), .B(G78gat), .ZN(new_n540));
  XOR2_X1   g339(.A(G57gat), .B(G64gat), .Z(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(KEYINPUT9), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT91), .B1(new_n547), .B2(new_n540), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550));
  INV_X1    g349(.A(G71gat), .ZN(new_n551));
  INV_X1    g350(.A(G78gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n550), .B(new_n546), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n541), .A2(new_n540), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n214), .B1(new_n559), .B2(new_n558), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n564), .A2(G183gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(G183gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n568), .B2(new_n572), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n396), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n568), .A2(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n569), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n563), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n577), .B1(new_n574), .B2(new_n575), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n573), .A3(new_n579), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n562), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n232), .A2(new_n234), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n592), .A3(KEYINPUT7), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n595), .A2(new_n602), .A3(new_n599), .A4(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n588), .A2(new_n606), .B1(KEYINPUT95), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n604), .A2(new_n605), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n230), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT41), .ZN(new_n612));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n609), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G134gat), .B(G162gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n608), .A2(KEYINPUT95), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n612), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n616), .B(new_n619), .Z(new_n620));
  NOR2_X1   g419(.A1(new_n587), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G230gat), .ZN(new_n622));
  INV_X1    g421(.A(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n544), .A2(new_n548), .B1(new_n556), .B2(new_n554), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n605), .A2(KEYINPUT96), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n606), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n625), .A3(new_n626), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT97), .B(KEYINPUT10), .Z(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n610), .A2(KEYINPUT98), .A3(KEYINPUT10), .A4(new_n625), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n558), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n624), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n622), .B(new_n623), .C1(new_n628), .C2(new_n629), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n354), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n639), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n539), .A2(new_n621), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n519), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n520), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n204), .A2(new_n207), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT42), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n652), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n649), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n652), .B2(KEYINPUT42), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n499), .A2(new_n501), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(G15gat), .B1(new_n646), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n537), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n646), .A2(G15gat), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n518), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n664), .B(new_n666), .ZN(G1327gat));
  NAND3_X1  g466(.A1(new_n587), .A2(new_n645), .A3(new_n258), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n616), .B(new_n619), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(KEYINPUT44), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n517), .A2(KEYINPUT102), .A3(new_n538), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT102), .B1(new_n517), .B2(new_n538), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n517), .A2(new_n538), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n620), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n668), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n352), .ZN(new_n679));
  INV_X1    g478(.A(new_n587), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n669), .A3(new_n644), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n539), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n219), .A3(new_n519), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n684), .ZN(G1328gat));
  OAI21_X1  g484(.A(G36gat), .B1(new_n678), .B2(new_n429), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n682), .A2(new_n220), .A3(new_n520), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n694));
  INV_X1    g493(.A(G43gat), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n677), .B2(new_n661), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n539), .A2(new_n681), .A3(new_n695), .A4(new_n659), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n693), .B(new_n694), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n668), .ZN(new_n701));
  INV_X1    g500(.A(new_n670), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n674), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n517), .A2(KEYINPUT102), .A3(new_n538), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n669), .B1(new_n517), .B2(new_n538), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n661), .B(new_n701), .C1(new_n706), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n697), .B(KEYINPUT104), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n711), .A2(new_n691), .A3(new_n692), .A4(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n700), .A2(new_n713), .ZN(G1330gat));
  AOI21_X1  g513(.A(G50gat), .B1(new_n682), .B2(new_n518), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n518), .A2(G50gat), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n677), .B2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g517(.A(new_n258), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n587), .A2(new_n620), .A3(new_n645), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n719), .B(new_n720), .C1(new_n671), .C2(new_n672), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n519), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n705), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n725), .A2(new_n719), .A3(new_n520), .A4(new_n720), .ZN(new_n726));
  NAND2_X1  g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT106), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n722), .A2(new_n730), .A3(new_n520), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n722), .A2(G71gat), .A3(new_n661), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n551), .B1(new_n721), .B2(new_n658), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n463), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n552), .ZN(G1335gat));
  OAI21_X1  g539(.A(KEYINPUT107), .B1(new_n680), .B2(new_n258), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n587), .A2(new_n742), .A3(new_n719), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n644), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n673), .B2(new_n676), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n352), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n707), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n744), .A2(new_n707), .A3(KEYINPUT51), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n644), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n519), .A2(new_n597), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n748), .B1(new_n755), .B2(new_n756), .ZN(G1336gat));
  NAND2_X1  g556(.A1(new_n746), .A2(new_n520), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n645), .A2(G92gat), .A3(new_n429), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n752), .B2(new_n754), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n751), .A2(new_n753), .B1(KEYINPUT108), .B2(new_n760), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n758), .A2(G92gat), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n747), .B2(new_n537), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n659), .A2(new_n473), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n755), .B2(new_n770), .ZN(G1338gat));
  NAND2_X1  g570(.A1(new_n746), .A2(new_n518), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n463), .A2(new_n645), .A3(G106gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n751), .A2(new_n753), .B1(KEYINPUT110), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n772), .A2(G106gat), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n772), .A2(G106gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n752), .B2(new_n754), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n777), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n780), .ZN(G1339gat));
  NAND2_X1  g580(.A1(new_n519), .A2(new_n429), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n631), .A2(new_n636), .A3(new_n624), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n637), .B2(KEYINPUT111), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n631), .A2(new_n636), .A3(new_n785), .A4(new_n624), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n637), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(new_n643), .ZN(new_n791));
  INV_X1    g590(.A(new_n643), .ZN(new_n792));
  AOI211_X1 g591(.A(KEYINPUT112), .B(new_n792), .C1(new_n637), .C2(new_n789), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n639), .A2(new_n643), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n787), .B(KEYINPUT55), .C1(new_n791), .C2(new_n793), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n258), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n245), .A2(new_n246), .A3(new_n244), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n240), .B1(new_n235), .B2(new_n239), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n253), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n803), .A2(new_n644), .A3(new_n257), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n669), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n803), .A2(new_n257), .A3(new_n804), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n620), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n587), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n621), .A2(new_n645), .A3(new_n719), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n782), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n463), .A2(new_n493), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n272), .A3(new_n258), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n518), .A2(new_n658), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n260), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1340gat));
  OAI21_X1  g625(.A(G120gat), .B1(new_n824), .B2(new_n645), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n644), .A2(new_n270), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT115), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n827), .B(new_n832), .C1(new_n820), .C2(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1341gat));
  NOR3_X1   g633(.A1(new_n824), .A2(new_n269), .A3(new_n587), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n821), .A2(new_n680), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n269), .B2(new_n836), .ZN(G1342gat));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n268), .A3(new_n620), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n824), .B2(new_n669), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n811), .A2(KEYINPUT117), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n796), .A2(new_n845), .A3(new_n797), .A4(new_n798), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n259), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n620), .B1(new_n847), .B2(new_n805), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n669), .A2(new_n812), .A3(new_n811), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n587), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n463), .B1(new_n850), .B2(new_n817), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n661), .A2(new_n782), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n680), .B1(new_n810), .B2(new_n814), .ZN(new_n855));
  NOR4_X1   g654(.A1(new_n587), .A2(new_n620), .A3(new_n644), .A4(new_n258), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n852), .B(new_n518), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n853), .A2(new_n258), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n843), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n518), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n260), .A2(G141gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT118), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n463), .B1(new_n816), .B2(new_n817), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n854), .A4(new_n862), .ZN(new_n867));
  INV_X1    g666(.A(new_n862), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n854), .B(new_n857), .C1(new_n851), .C2(new_n852), .ZN(new_n871));
  OAI21_X1  g670(.A(G141gat), .B1(new_n871), .B2(new_n260), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n859), .A2(new_n864), .B1(new_n873), .B2(new_n843), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n861), .A2(new_n286), .A3(new_n644), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n621), .A2(new_n645), .A3(new_n260), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n850), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n518), .B1(new_n855), .B2(new_n856), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n878), .A2(new_n518), .B1(new_n879), .B2(KEYINPUT57), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n854), .B(KEYINPUT120), .Z(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n644), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n876), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n876), .B(G148gat), .C1(new_n871), .C2(new_n645), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n875), .B1(new_n883), .B2(new_n885), .ZN(G1345gat));
  XNOR2_X1  g685(.A(KEYINPUT72), .B(G155gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n680), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT122), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n861), .A2(new_n680), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT121), .ZN(new_n892));
  INV_X1    g691(.A(new_n887), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1346gat));
  AOI21_X1  g693(.A(G162gat), .B1(new_n861), .B2(new_n620), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n871), .A2(new_n669), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n519), .A2(new_n429), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n823), .B(new_n898), .C1(new_n855), .C2(new_n856), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n260), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n819), .A2(KEYINPUT123), .A3(new_n520), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT123), .B1(new_n819), .B2(new_n520), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n519), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(new_n903), .C1(new_n855), .C2(new_n856), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n258), .A2(new_n384), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT124), .ZN(G1348gat));
  NOR3_X1   g706(.A1(new_n899), .A2(new_n354), .A3(new_n645), .ZN(new_n908));
  INV_X1    g707(.A(new_n904), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n644), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n354), .B2(new_n910), .ZN(G1349gat));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n680), .A2(new_n375), .ZN(new_n913));
  OR3_X1    g712(.A1(new_n904), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n904), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G183gat), .B1(new_n899), .B2(new_n587), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT60), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n909), .A2(new_n376), .A3(new_n620), .ZN(new_n923));
  OAI21_X1  g722(.A(G190gat), .B1(new_n899), .B2(new_n669), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  NAND2_X1  g727(.A1(new_n898), .A2(new_n537), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n880), .A2(new_n259), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G197gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n865), .A2(new_n930), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n933), .A2(G197gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n719), .B2(new_n934), .ZN(G1352gat));
  OR3_X1    g734(.A1(new_n933), .A2(G204gat), .A3(new_n645), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT126), .B1(new_n936), .B2(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n880), .A2(new_n644), .A3(new_n930), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G204gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n933), .A2(G204gat), .A3(new_n645), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n937), .A2(new_n938), .A3(new_n940), .A4(new_n944), .ZN(G1353gat));
  OR3_X1    g744(.A1(new_n933), .A2(new_n587), .A3(new_n408), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n880), .A2(new_n680), .A3(new_n930), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  NAND2_X1  g749(.A1(new_n878), .A2(new_n518), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n879), .A2(KEYINPUT57), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n930), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n620), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n953), .B1(new_n880), .B2(new_n930), .ZN(new_n956));
  OAI21_X1  g755(.A(G218gat), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n620), .A2(new_n394), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n933), .B2(new_n958), .ZN(G1355gat));
endmodule


