

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  NOR2_X1 U322 ( .A1(n580), .A2(n486), .ZN(n487) );
  XNOR2_X1 U323 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U324 ( .A(KEYINPUT28), .B(n467), .Z(n529) );
  INV_X1 U325 ( .A(KEYINPUT46), .ZN(n362) );
  XNOR2_X1 U326 ( .A(n362), .B(KEYINPUT114), .ZN(n363) );
  XNOR2_X1 U327 ( .A(n364), .B(n363), .ZN(n381) );
  INV_X1 U328 ( .A(KEYINPUT86), .ZN(n298) );
  XNOR2_X1 U329 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U330 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U331 ( .A(n335), .B(n334), .ZN(n336) );
  NOR2_X1 U332 ( .A1(n531), .A2(n452), .ZN(n560) );
  XNOR2_X1 U333 ( .A(n341), .B(n398), .ZN(n570) );
  XNOR2_X1 U334 ( .A(n429), .B(n308), .ZN(n531) );
  XNOR2_X1 U335 ( .A(n490), .B(n489), .ZN(n501) );
  XNOR2_X1 U336 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U337 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT0), .B(G134GAT), .Z(n291) );
  XNOR2_X1 U339 ( .A(KEYINPUT84), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(n292), .ZN(n429) );
  XOR2_X1 U342 ( .A(G176GAT), .B(KEYINPUT87), .Z(n294) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U345 ( .A(G120GAT), .B(G71GAT), .Z(n359) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(G99GAT), .Z(n296) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G190GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U349 ( .A(n359), .B(n297), .Z(n301) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U351 ( .A(G183GAT), .B(KEYINPUT18), .Z(n303) );
  XNOR2_X1 U352 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n316) );
  XNOR2_X1 U354 ( .A(n316), .B(KEYINPUT85), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U356 ( .A(n307), .B(n306), .Z(n308) );
  XOR2_X1 U357 ( .A(G169GAT), .B(G8GAT), .Z(n329) );
  XOR2_X1 U358 ( .A(G176GAT), .B(G64GAT), .Z(n351) );
  XNOR2_X1 U359 ( .A(n329), .B(n351), .ZN(n320) );
  XOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .Z(n385) );
  XOR2_X1 U361 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n310) );
  XNOR2_X1 U362 ( .A(G204GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U364 ( .A(n385), .B(n311), .Z(n313) );
  NAND2_X1 U365 ( .A1(G226GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U367 ( .A(G211GAT), .B(KEYINPUT21), .Z(n315) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n443) );
  XOR2_X1 U370 ( .A(n316), .B(n443), .Z(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n519) );
  XOR2_X1 U373 ( .A(G22GAT), .B(G141GAT), .Z(n322) );
  XNOR2_X1 U374 ( .A(G50GAT), .B(G36GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U376 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n324) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(G113GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U379 ( .A(n326), .B(n325), .Z(n337) );
  XOR2_X1 U380 ( .A(G1GAT), .B(KEYINPUT70), .Z(n328) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(KEYINPUT71), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n369) );
  XOR2_X1 U383 ( .A(n329), .B(n369), .Z(n335) );
  XOR2_X1 U384 ( .A(KEYINPUT30), .B(KEYINPUT72), .Z(n331) );
  XNOR2_X1 U385 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n333) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U389 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n339) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(KEYINPUT7), .B(n340), .ZN(n398) );
  INV_X1 U393 ( .A(n570), .ZN(n457) );
  XOR2_X1 U394 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n343) );
  NAND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(n344), .B(KEYINPUT75), .Z(n350) );
  XOR2_X1 U398 ( .A(G78GAT), .B(G148GAT), .Z(n346) );
  XNOR2_X1 U399 ( .A(G106GAT), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n445) );
  XOR2_X1 U401 ( .A(KEYINPUT76), .B(G92GAT), .Z(n348) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n393) );
  XNOR2_X1 U404 ( .A(n445), .B(n393), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT79), .B(KEYINPUT74), .Z(n353) );
  XOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .Z(n367) );
  XNOR2_X1 U408 ( .A(n351), .B(n367), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U411 ( .A(KEYINPUT31), .B(KEYINPUT78), .Z(n357) );
  XNOR2_X1 U412 ( .A(KEYINPUT77), .B(KEYINPUT73), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n573) );
  XNOR2_X1 U416 ( .A(n573), .B(KEYINPUT41), .ZN(n504) );
  NOR2_X1 U417 ( .A1(n457), .A2(n504), .ZN(n364) );
  XOR2_X1 U418 ( .A(KEYINPUT14), .B(G64GAT), .Z(n366) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(G183GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U421 ( .A(n368), .B(n367), .Z(n371) );
  XOR2_X1 U422 ( .A(G22GAT), .B(G155GAT), .Z(n437) );
  XNOR2_X1 U423 ( .A(n369), .B(n437), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U425 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n373) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U428 ( .A(n375), .B(n374), .Z(n380) );
  XOR2_X1 U429 ( .A(G211GAT), .B(G78GAT), .Z(n377) );
  XNOR2_X1 U430 ( .A(G127GAT), .B(G71GAT), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n378), .B(KEYINPUT15), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n484) );
  NAND2_X1 U434 ( .A1(n381), .A2(n484), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n382), .B(KEYINPUT115), .ZN(n400) );
  XOR2_X1 U436 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n384) );
  XNOR2_X1 U437 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n386) );
  XOR2_X1 U439 ( .A(n386), .B(n385), .Z(n388) );
  XNOR2_X1 U440 ( .A(G134GAT), .B(G106GAT), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n397) );
  XOR2_X1 U442 ( .A(KEYINPUT82), .B(KEYINPUT9), .Z(n390) );
  NAND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U445 ( .A(n391), .B(KEYINPUT81), .Z(n395) );
  XNOR2_X1 U446 ( .A(G50GAT), .B(KEYINPUT80), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n392), .B(G162GAT), .ZN(n440) );
  XNOR2_X1 U448 ( .A(n440), .B(n393), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n399) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n540) );
  NAND2_X1 U452 ( .A1(n400), .A2(n540), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n401), .B(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U454 ( .A(KEYINPUT36), .B(n540), .ZN(n580) );
  NOR2_X1 U455 ( .A1(n484), .A2(n580), .ZN(n403) );
  XOR2_X1 U456 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  NAND2_X1 U458 ( .A1(n457), .A2(n404), .ZN(n405) );
  NOR2_X1 U459 ( .A1(n405), .A2(n573), .ZN(n406) );
  NOR2_X1 U460 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U461 ( .A(KEYINPUT48), .B(n408), .ZN(n528) );
  NOR2_X1 U462 ( .A1(n519), .A2(n528), .ZN(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT54), .B(n409), .ZN(n433) );
  XOR2_X1 U464 ( .A(KEYINPUT95), .B(KEYINPUT98), .Z(n411) );
  XNOR2_X1 U465 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U467 ( .A(G57GAT), .B(G155GAT), .Z(n413) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G120GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n423) );
  XOR2_X1 U471 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n417) );
  XNOR2_X1 U472 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(G141GAT), .B(n418), .Z(n446) );
  XOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT4), .B(KEYINPUT97), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n446), .B(n421), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n432) );
  XOR2_X1 U480 ( .A(G85GAT), .B(G162GAT), .Z(n425) );
  XNOR2_X1 U481 ( .A(G29GAT), .B(G148GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT1), .B(n426), .Z(n428) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U486 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n517) );
  NAND2_X1 U488 ( .A1(n433), .A2(n517), .ZN(n568) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n435) );
  XNOR2_X1 U490 ( .A(KEYINPUT89), .B(KEYINPUT93), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U492 ( .A(n436), .B(KEYINPUT22), .Z(n439) );
  XNOR2_X1 U493 ( .A(n437), .B(KEYINPUT88), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n450) );
  XOR2_X1 U495 ( .A(KEYINPUT90), .B(n440), .Z(n442) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n467) );
  NOR2_X1 U502 ( .A1(n568), .A2(n467), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  INV_X1 U504 ( .A(n504), .ZN(n548) );
  NAND2_X1 U505 ( .A1(n560), .A2(n548), .ZN(n456) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n453) );
  NOR2_X1 U508 ( .A1(n573), .A2(n457), .ZN(n488) );
  XOR2_X1 U509 ( .A(KEYINPUT27), .B(n519), .Z(n466) );
  XOR2_X1 U510 ( .A(KEYINPUT26), .B(KEYINPUT101), .Z(n459) );
  NAND2_X1 U511 ( .A1(n531), .A2(n467), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n567) );
  INV_X1 U513 ( .A(n567), .ZN(n545) );
  NAND2_X1 U514 ( .A1(n466), .A2(n545), .ZN(n464) );
  XNOR2_X1 U515 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n531), .A2(n519), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n467), .A2(n460), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n465), .A2(n517), .ZN(n470) );
  INV_X1 U521 ( .A(n531), .ZN(n496) );
  INV_X1 U522 ( .A(n517), .ZN(n491) );
  NAND2_X1 U523 ( .A1(n491), .A2(n466), .ZN(n527) );
  NOR2_X1 U524 ( .A1(n496), .A2(n527), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n468), .A2(n529), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n470), .A2(n469), .ZN(n483) );
  INV_X1 U527 ( .A(n484), .ZN(n576) );
  NAND2_X1 U528 ( .A1(n540), .A2(n576), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  AND2_X1 U530 ( .A1(n483), .A2(n472), .ZN(n505) );
  NAND2_X1 U531 ( .A1(n488), .A2(n505), .ZN(n479) );
  NOR2_X1 U532 ( .A1(n517), .A2(n479), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT34), .B(n473), .Z(n474) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n519), .A2(n479), .ZN(n475) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n475), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n531), .A2(n479), .ZN(n477) );
  XNOR2_X1 U538 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U540 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NOR2_X1 U541 ( .A1(n529), .A2(n479), .ZN(n480) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n480), .Z(G1327GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT104), .B(KEYINPUT107), .Z(n482) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(n493) );
  XOR2_X1 U546 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n490) );
  NAND2_X1 U547 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U548 ( .A(KEYINPUT105), .B(n485), .Z(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n487), .Z(n516) );
  NAND2_X1 U550 ( .A1(n488), .A2(n516), .ZN(n489) );
  NAND2_X1 U551 ( .A1(n491), .A2(n501), .ZN(n492) );
  XOR2_X1 U552 ( .A(n493), .B(n492), .Z(G1328GAT) );
  INV_X1 U553 ( .A(n519), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n494), .A2(n501), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n498) );
  NAND2_X1 U557 ( .A1(n501), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U559 ( .A(n499), .B(G43GAT), .Z(G1330GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT109), .Z(n503) );
  INV_X1 U561 ( .A(n529), .ZN(n500) );
  NAND2_X1 U562 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n570), .A2(n504), .ZN(n515) );
  NAND2_X1 U565 ( .A1(n515), .A2(n505), .ZN(n512) );
  NOR2_X1 U566 ( .A1(n517), .A2(n512), .ZN(n507) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NOR2_X1 U570 ( .A1(n519), .A2(n512), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n531), .A2(n512), .ZN(n511) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n529), .A2(n512), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n523) );
  NOR2_X1 U579 ( .A1(n517), .A2(n523), .ZN(n518) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n531), .A2(n523), .ZN(n521) );
  XOR2_X1 U584 ( .A(KEYINPUT112), .B(n521), .Z(n522) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n523), .ZN(n525) );
  XNOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n544), .A2(n529), .ZN(n530) );
  NOR2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U593 ( .A(KEYINPUT116), .B(n532), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n541), .A2(n570), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U597 ( .A1(n548), .A2(n541), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n537) );
  NAND2_X1 U601 ( .A1(n541), .A2(n576), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  INV_X1 U605 ( .A(n540), .ZN(n559) );
  NAND2_X1 U606 ( .A1(n559), .A2(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT119), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n554), .A2(n570), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n550) );
  NAND2_X1 U614 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n576), .A2(n554), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT121), .Z(n556) );
  NAND2_X1 U620 ( .A1(n554), .A2(n559), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n560), .A2(n570), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n576), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n565) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(n566), .Z(n572) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT124), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n570), .A2(n578), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n578), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n578), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n582) );
  INV_X1 U644 ( .A(n578), .ZN(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

