//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT90), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT0), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(KEYINPUT0), .B2(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G146), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n197), .A2(KEYINPUT65), .A3(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n204), .A3(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n196), .A2(new_n203), .B1(new_n206), .B2(KEYINPUT0), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n198), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G128), .A3(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n203), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT68), .B1(new_n216), .B2(new_n203), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n208), .B(new_n211), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n209), .B1(new_n219), .B2(KEYINPUT86), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n203), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n216), .A2(KEYINPUT68), .A3(new_n203), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n210), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n208), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G224), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT7), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n209), .B2(KEYINPUT89), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT2), .B(G113), .Z(new_n235));
  XNOR2_X1  g049(.A(G116), .B(G119), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT69), .B1(new_n235), .B2(new_n236), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n240));
  INV_X1    g054(.A(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G104), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G107), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n240), .A2(new_n247), .A3(new_n241), .A4(G104), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n243), .A2(new_n244), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n246), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(G107), .ZN(new_n251));
  OAI21_X1  g065(.A(G101), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  OR3_X1    g069(.A1(new_n255), .A2(KEYINPUT5), .A3(G119), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(G113), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n239), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G122), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT8), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n237), .A2(new_n238), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n236), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(G113), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n254), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n261), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n258), .B(new_n260), .C1(new_n253), .C2(new_n266), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n237), .A2(new_n238), .B1(new_n235), .B2(new_n236), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n248), .A2(new_n246), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n247), .B1(new_n251), .B2(new_n240), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT80), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n243), .A2(new_n273), .A3(new_n246), .A4(new_n248), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n272), .A3(G101), .A4(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(G101), .A3(new_n274), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n277), .A2(KEYINPUT81), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT81), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n253), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n239), .A2(new_n282), .A3(new_n257), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n283), .A3(new_n259), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n220), .A2(new_n227), .A3(new_n232), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n234), .A2(new_n267), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n220), .A2(new_n230), .A3(new_n227), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n230), .B1(new_n220), .B2(new_n227), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT85), .A2(KEYINPUT6), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n259), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n268), .A2(new_n275), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n277), .A2(new_n278), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n277), .A2(KEYINPUT81), .A3(new_n278), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n283), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n259), .B1(new_n281), .B2(new_n283), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n293), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n291), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT87), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n288), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n289), .A2(new_n290), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n284), .B2(new_n293), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n303), .A2(new_n292), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT87), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n188), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n286), .A2(new_n287), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n313), .B2(KEYINPUT87), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n306), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n308), .A3(new_n310), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n187), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G478), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT15), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n190), .A2(KEYINPUT13), .A3(G143), .ZN(new_n325));
  INV_X1    g139(.A(G134), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G128), .B(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n326), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT97), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n327), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n331), .B2(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT96), .B1(new_n255), .B2(G122), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT96), .ZN(new_n335));
  INV_X1    g149(.A(G122), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G116), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n255), .A2(G122), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G107), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n241), .A3(new_n339), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT9), .B(G234), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n345), .A2(new_n346), .A3(G953), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n338), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT98), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n338), .A2(KEYINPUT98), .A3(new_n348), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n351), .B(new_n352), .C1(KEYINPUT14), .C2(new_n339), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(G107), .ZN(new_n354));
  INV_X1    g168(.A(new_n330), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n328), .A2(new_n326), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n342), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n344), .B(new_n347), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n347), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n353), .B2(G107), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n333), .A2(new_n343), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n324), .B1(new_n363), .B2(new_n287), .ZN(new_n364));
  AOI211_X1 g178(.A(G902), .B(new_n323), .C1(new_n358), .C2(new_n362), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n208), .A2(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT16), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(G146), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(G146), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n375));
  INV_X1    g189(.A(G131), .ZN(new_n376));
  NOR2_X1   g190(.A1(G237), .A2(G953), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G214), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n200), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT91), .A2(G143), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT91), .A2(G143), .ZN(new_n382));
  OAI211_X1 g196(.A(G214), .B(new_n377), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n376), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT17), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n374), .B(new_n375), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n371), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n197), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n370), .A2(new_n371), .A3(G146), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI211_X1 g205(.A(new_n386), .B(new_n376), .C1(new_n380), .C2(new_n383), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT94), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n380), .A2(new_n383), .A3(new_n376), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n387), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n380), .A2(new_n383), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n397), .A2(KEYINPUT18), .A3(G131), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(KEYINPUT18), .B2(G131), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n368), .A2(new_n369), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G146), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n368), .A2(new_n369), .A3(new_n197), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OR3_X1    g217(.A1(new_n398), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT93), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(new_n245), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n400), .B(KEYINPUT19), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n390), .B1(new_n410), .B2(G146), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT92), .ZN(new_n412));
  INV_X1    g226(.A(new_n394), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n384), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n385), .A2(KEYINPUT92), .A3(new_n394), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n398), .A2(new_n399), .A3(new_n403), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n409), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n408), .A2(new_n418), .A3(KEYINPUT95), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n421), .A2(KEYINPUT20), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n422), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n408), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n407), .B1(new_n396), .B2(new_n404), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n287), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G475), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n366), .A2(new_n424), .A3(new_n427), .A4(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(KEYINPUT99), .A2(G952), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT99), .A2(G952), .ZN(new_n435));
  AOI21_X1  g249(.A(G953), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G234), .ZN(new_n437));
  INV_X1    g251(.A(G237), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(G898), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n287), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT100), .B1(new_n432), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n424), .A2(new_n427), .A3(new_n431), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT100), .ZN(new_n446));
  INV_X1    g260(.A(new_n443), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n366), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n321), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G472), .A2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT66), .A2(G137), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(KEYINPUT66), .A2(G137), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT11), .ZN(new_n461));
  NOR4_X1   g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n326), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n326), .B2(G137), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n326), .A2(G137), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G131), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n460), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(KEYINPUT11), .A3(G134), .A4(new_n458), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(new_n376), .A3(new_n463), .A4(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n457), .B1(new_n470), .B2(new_n207), .ZN(new_n471));
  AOI21_X1  g285(.A(G134), .B1(new_n467), .B2(new_n458), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n326), .A2(G137), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n225), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n198), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n199), .A2(new_n200), .A3(G146), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n480), .A2(new_n195), .B1(new_n189), .B2(new_n205), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n469), .B2(new_n466), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n211), .B1(new_n217), .B2(new_n218), .ZN(new_n483));
  INV_X1    g297(.A(new_n475), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n476), .B(new_n268), .C1(new_n485), .C2(KEYINPUT30), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT26), .B(G101), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n377), .A2(G210), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n268), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT71), .B1(new_n486), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT31), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n486), .A2(new_n494), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT31), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n485), .A2(new_n493), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n268), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n485), .A2(new_n493), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n491), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n456), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  AOI211_X1 g325(.A(KEYINPUT73), .B(new_n509), .C1(new_n497), .C2(new_n500), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n455), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n491), .A3(new_n508), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n486), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n492), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n508), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n503), .A2(new_n504), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(KEYINPUT28), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n492), .A2(new_n515), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n287), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G472), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n498), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n494), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n499), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n500), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n510), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n501), .A2(new_n456), .A3(new_n510), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n453), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n513), .B(new_n525), .C1(new_n534), .C2(KEYINPUT32), .ZN(new_n535));
  OAI21_X1  g349(.A(G221), .B1(new_n345), .B2(G902), .ZN(new_n536));
  INV_X1    g350(.A(G469), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n282), .A2(KEYINPUT10), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n190), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n198), .A2(new_n204), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n211), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n282), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n543));
  AOI22_X1  g357(.A1(new_n538), .A2(new_n483), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n470), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n279), .A2(new_n280), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n275), .A2(new_n207), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n211), .B(new_n253), .C1(new_n217), .C2(new_n218), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n542), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n545), .B2(KEYINPUT83), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n550), .A2(new_n470), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n550), .B2(new_n470), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G140), .ZN(new_n556));
  INV_X1    g370(.A(G227), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n538), .A2(new_n483), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n542), .A2(new_n543), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n547), .B1(new_n299), .B2(new_n300), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n470), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n559), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n548), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n537), .B1(new_n568), .B2(new_n287), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n548), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n559), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n548), .B(new_n566), .C1(new_n553), .C2(new_n554), .ZN(new_n572));
  AOI211_X1 g386(.A(G469), .B(G902), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n536), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n536), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n548), .A2(new_n566), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n565), .A2(new_n578), .B1(new_n555), .B2(new_n559), .ZN(new_n579));
  OAI21_X1  g393(.A(G469), .B1(new_n579), .B2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n572), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n537), .A3(new_n287), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT84), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT22), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G137), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n190), .A2(G119), .ZN(new_n590));
  INV_X1    g404(.A(G119), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G128), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT74), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(KEYINPUT23), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(KEYINPUT23), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT23), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT74), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n595), .A2(new_n597), .A3(G119), .A4(new_n190), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n598), .A3(G110), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n590), .A2(new_n592), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT24), .B(G110), .Z(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n589), .B1(new_n374), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n599), .A2(new_n602), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n391), .A3(KEYINPUT75), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n594), .A2(new_n598), .ZN(new_n607));
  OAI22_X1  g421(.A1(new_n607), .A2(G110), .B1(new_n600), .B2(new_n601), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n390), .A2(new_n402), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n604), .A2(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n588), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n604), .A2(new_n606), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(KEYINPUT76), .A3(new_n588), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n346), .B1(G234), .B2(new_n287), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT78), .Z(new_n623));
  INV_X1    g437(.A(KEYINPUT77), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n617), .B2(new_n618), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT25), .B(G902), .C1(new_n617), .C2(new_n618), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n619), .A2(new_n287), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT25), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n625), .A2(new_n626), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(KEYINPUT77), .A3(new_n632), .A4(new_n620), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n623), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n451), .A2(new_n535), .A3(new_n585), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  NAND2_X1  g451(.A1(new_n313), .A2(KEYINPUT87), .ZN(new_n638));
  AND4_X1   g452(.A1(new_n187), .A2(new_n638), .A3(new_n319), .A4(new_n288), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n187), .B1(new_n317), .B2(new_n319), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n450), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT101), .ZN(new_n642));
  AOI21_X1  g456(.A(G478), .B1(new_n363), .B2(new_n287), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n358), .A2(KEYINPUT33), .A3(new_n362), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT33), .B1(new_n358), .B2(new_n362), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n322), .A2(G902), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n445), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n450), .C1(new_n639), .C2(new_n640), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n642), .A2(new_n447), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n287), .B1(new_n511), .B2(new_n512), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n532), .A2(new_n533), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n654), .A2(G472), .B1(new_n655), .B2(new_n452), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n656), .A2(new_n585), .A3(new_n635), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G6));
  AND2_X1   g475(.A1(new_n424), .A2(new_n431), .ZN(new_n662));
  INV_X1    g476(.A(new_n366), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n421), .A2(new_n423), .ZN(new_n664));
  INV_X1    g478(.A(new_n422), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n426), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n642), .A2(new_n447), .A3(new_n651), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n657), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT35), .B(G107), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT103), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n670), .B(new_n672), .ZN(G9));
  INV_X1    g487(.A(KEYINPUT36), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n588), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n610), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n621), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n629), .A2(new_n633), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n451), .A2(new_n656), .A3(new_n585), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(new_n187), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n309), .B2(new_n314), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n320), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n650), .B1(new_n684), .B2(new_n450), .ZN(new_n685));
  INV_X1    g499(.A(new_n450), .ZN(new_n686));
  AOI211_X1 g500(.A(KEYINPUT101), .B(new_n686), .C1(new_n683), .C2(new_n320), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n629), .A2(new_n633), .A3(new_n677), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n655), .A2(new_n455), .B1(G472), .B2(new_n524), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n452), .B1(new_n511), .B2(new_n512), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n454), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n439), .B(KEYINPUT105), .Z(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(G900), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(G900), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n442), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT106), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n667), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n688), .A2(new_n693), .A3(new_n585), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XOR2_X1   g517(.A(new_n700), .B(KEYINPUT107), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT39), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n585), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT108), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n321), .B(KEYINPUT38), .Z(new_n714));
  AOI21_X1  g528(.A(KEYINPUT32), .B1(new_n655), .B2(new_n452), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n495), .A2(new_n496), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n520), .A2(new_n492), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n287), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G472), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n513), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n424), .A2(new_n427), .A3(new_n431), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n663), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n689), .A2(new_n450), .A3(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n714), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n711), .A2(new_n713), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  INV_X1    g543(.A(new_n649), .ZN(new_n730));
  INV_X1    g544(.A(new_n700), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n688), .A2(new_n693), .A3(new_n585), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  NAND2_X1  g548(.A1(new_n581), .A2(new_n287), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n536), .A3(new_n582), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n513), .A2(new_n525), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n635), .B(new_n738), .C1(new_n715), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n652), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT110), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n741), .B(new_n743), .ZN(G15));
  NOR2_X1   g558(.A1(new_n668), .A2(new_n740), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n255), .ZN(G18));
  NAND3_X1  g560(.A1(new_n535), .A2(new_n449), .A3(new_n678), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n642), .A2(new_n651), .A3(new_n738), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n591), .ZN(G21));
  NAND3_X1  g564(.A1(new_n642), .A2(new_n651), .A3(new_n725), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n521), .A2(new_n491), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n453), .B1(new_n752), .B2(new_n501), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n654), .B2(G472), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n737), .A2(new_n443), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n635), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n336), .ZN(G24));
  AOI211_X1 g572(.A(new_n753), .B(new_n689), .C1(G472), .C2(new_n654), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n688), .A2(new_n759), .A3(new_n732), .A4(new_n738), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT111), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  AND4_X1   g576(.A1(new_n450), .A2(new_n583), .A3(new_n315), .A4(new_n320), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n535), .A2(new_n635), .A3(new_n732), .A4(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n634), .B1(new_n690), .B2(new_n692), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(KEYINPUT42), .A3(new_n732), .A4(new_n763), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n376), .ZN(G33));
  NAND4_X1  g588(.A1(new_n535), .A2(new_n635), .A3(new_n701), .A4(new_n763), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  NAND2_X1  g590(.A1(new_n579), .A2(KEYINPUT45), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT113), .ZN(new_n778));
  OAI21_X1  g592(.A(G469), .B1(new_n579), .B2(KEYINPUT45), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(KEYINPUT113), .B2(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(G469), .A2(G902), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n573), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n782), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(new_n536), .A3(new_n705), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n321), .A2(new_n686), .ZN(new_n788));
  INV_X1    g602(.A(new_n656), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n723), .A2(new_n648), .B1(KEYINPUT114), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n643), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n644), .A2(new_n645), .ZN(new_n793));
  INV_X1    g607(.A(new_n647), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n445), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT114), .B(KEYINPUT43), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(new_n678), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT44), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(KEYINPUT44), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n787), .A2(new_n788), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NAND2_X1  g618(.A1(new_n786), .A2(new_n536), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n786), .A2(new_n807), .A3(new_n536), .ZN(new_n808));
  INV_X1    g622(.A(new_n788), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n732), .A2(new_n634), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n535), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  NOR3_X1   g627(.A1(new_n796), .A2(new_n686), .A3(new_n577), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n736), .A2(new_n582), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n635), .B(new_n814), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT115), .Z(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n714), .A3(new_n722), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n678), .A2(new_n574), .A3(new_n731), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n715), .B2(new_n721), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n751), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n689), .A2(new_n583), .A3(new_n700), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n655), .A2(new_n455), .B1(G472), .B2(new_n719), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n692), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n688), .A3(new_n829), .A4(new_n725), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n702), .A2(new_n760), .A3(new_n733), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n825), .A2(new_n830), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n535), .A2(new_n585), .A3(new_n678), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n688), .C1(new_n701), .C2(new_n732), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT52), .A4(new_n760), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n747), .A2(new_n748), .B1(new_n751), .B2(new_n756), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n741), .A3(new_n745), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n662), .A2(new_n366), .A3(new_n666), .A4(new_n700), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n576), .B2(new_n584), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n730), .A2(new_n574), .A3(new_n731), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n535), .A2(new_n843), .B1(new_n754), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n788), .A2(new_n678), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n775), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n723), .A2(new_n648), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n447), .A3(new_n432), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n686), .B(new_n849), .C1(new_n315), .C2(new_n320), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n656), .A3(new_n585), .A4(new_n635), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n636), .A2(new_n851), .A3(new_n679), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n841), .A2(new_n771), .A3(new_n853), .A4(new_n772), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n838), .A2(new_n839), .A3(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n771), .A2(new_n841), .A3(new_n772), .A4(new_n853), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n833), .A2(new_n837), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n839), .B1(new_n838), .B2(new_n854), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n839), .B1(new_n766), .B2(new_n768), .ZN(new_n861));
  INV_X1    g675(.A(new_n741), .ZN(new_n862));
  INV_X1    g676(.A(new_n745), .ZN(new_n863));
  INV_X1    g677(.A(new_n747), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n685), .A2(new_n687), .A3(new_n737), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n685), .A2(new_n687), .A3(new_n724), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n654), .A2(G472), .ZN(new_n867));
  INV_X1    g681(.A(new_n753), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n635), .A2(new_n867), .A3(new_n868), .A4(new_n755), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n864), .A2(new_n865), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n847), .B2(new_n852), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT54), .B1(new_n875), .B2(new_n857), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n860), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n859), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  INV_X1    g693(.A(new_n694), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n798), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT118), .Z(new_n882));
  AND2_X1   g696(.A1(new_n754), .A2(new_n635), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n714), .A2(new_n686), .A3(new_n738), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT119), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n886), .B(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n809), .A2(new_n737), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n634), .A2(new_n439), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n722), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n445), .A3(new_n648), .ZN(new_n894));
  INV_X1    g708(.A(new_n759), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n882), .A2(new_n890), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n889), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n806), .A2(new_n808), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n815), .A2(new_n536), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n809), .B(new_n884), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n879), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n884), .A2(new_n748), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT120), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n882), .A2(new_n767), .A3(new_n890), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT48), .Z(new_n906));
  OAI21_X1  g720(.A(new_n436), .B1(new_n892), .B2(new_n730), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n897), .A2(new_n901), .A3(new_n879), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n878), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n821), .B1(new_n911), .B2(new_n912), .ZN(G75));
  NAND2_X1  g727(.A1(new_n875), .A2(new_n857), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n860), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(G902), .A3(new_n188), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n318), .B(new_n310), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT56), .B1(new_n919), .B2(KEYINPUT121), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n229), .A2(G952), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n915), .A2(G902), .ZN(new_n927));
  INV_X1    g741(.A(G210), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n918), .B2(new_n929), .ZN(G51));
  INV_X1    g744(.A(new_n924), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n535), .A2(new_n843), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n754), .A2(new_n844), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n846), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n775), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n636), .A2(new_n851), .A3(new_n679), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT117), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n847), .A2(new_n852), .A3(new_n872), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n841), .B(new_n861), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n933), .B1(new_n838), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n932), .B1(new_n943), .B2(new_n858), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n838), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n945), .B2(new_n858), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n860), .A2(new_n876), .A3(KEYINPUT123), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n782), .B(KEYINPUT57), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n581), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n927), .A2(new_n781), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n931), .B1(new_n951), .B2(new_n952), .ZN(G54));
  NAND4_X1  g767(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n664), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n924), .B1(new_n954), .B2(new_n664), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n954), .B2(new_n664), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G60));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n859), .B2(new_n877), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n924), .B1(new_n962), .B2(new_n646), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n793), .A2(new_n961), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n948), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT60), .Z(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n945), .B2(new_n858), .ZN(new_n969));
  INV_X1    g783(.A(new_n619), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n931), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n676), .B(new_n968), .C1(new_n945), .C2(new_n858), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(KEYINPUT61), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n915), .A2(new_n974), .A3(new_n676), .A4(new_n968), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(G66));
  NAND2_X1  g793(.A1(new_n841), .A2(new_n939), .ZN(new_n980));
  NAND2_X1  g794(.A1(G224), .A2(G953), .ZN(new_n981));
  OAI22_X1  g795(.A1(new_n980), .A2(G953), .B1(new_n441), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n304), .B(new_n306), .C1(G898), .C2(new_n229), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G69));
  NAND3_X1  g798(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n985));
  INV_X1    g799(.A(new_n476), .ZN(new_n986));
  INV_X1    g800(.A(new_n485), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n457), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(new_n410), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n832), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n728), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n728), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n848), .A2(new_n432), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n707), .A2(new_n767), .A3(new_n788), .A4(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n803), .A2(new_n812), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n993), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n985), .B(new_n990), .C1(new_n999), .C2(G953), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n557), .A2(G900), .A3(G953), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n787), .A2(new_n767), .A3(new_n866), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n803), .A2(new_n812), .A3(new_n775), .A4(new_n1002), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1003), .A2(new_n773), .A3(new_n832), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n989), .B(new_n1001), .C1(new_n1004), .C2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1000), .A2(new_n1005), .ZN(G72));
  XOR2_X1   g820(.A(new_n516), .B(KEYINPUT127), .Z(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n491), .ZN(new_n1008));
  INV_X1    g822(.A(new_n980), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n993), .A2(new_n1009), .A3(new_n995), .A4(new_n998), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1012), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n1007), .A2(new_n491), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n924), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n855), .A2(new_n858), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n716), .A2(new_n517), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1018), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1013), .A2(new_n1017), .A3(new_n1020), .ZN(G57));
endmodule


