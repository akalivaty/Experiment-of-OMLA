//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n208), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NOR2_X1   g0042(.A1(G20), .A2(G33), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  AOI22_X1  g0044(.A1(new_n243), .A2(G50), .B1(G20), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT64), .B(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n245), .B1(new_n247), .B2(new_n202), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT11), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n248), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n255));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(new_n209), .A3(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n244), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n257), .A2(new_n251), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G68), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n254), .A2(new_n255), .A3(new_n259), .A4(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT14), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT13), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n214), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n214), .A2(new_n268), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G238), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT70), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT66), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n250), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n214), .A2(KEYINPUT66), .A3(new_n268), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n227), .A2(G1698), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G226), .B2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G97), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n283), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n266), .B1(new_n277), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n275), .A2(new_n276), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT70), .B1(new_n272), .B2(new_n274), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n294), .B(new_n266), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n265), .B(G169), .C1(new_n295), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT13), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G179), .A3(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n298), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n265), .B1(new_n305), .B2(G169), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n264), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n264), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n302), .B2(new_n298), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT3), .B(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G222), .A2(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G1698), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G223), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n283), .B(new_n320), .C1(G77), .C2(new_n316), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n279), .A2(new_n250), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n322), .A2(new_n267), .A3(new_n270), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n271), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(G226), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G190), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n243), .A2(G150), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n329), .B1(new_n209), .B2(new_n201), .C1(new_n247), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n251), .ZN(new_n332));
  INV_X1    g0132(.A(G50), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n261), .B2(G20), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n260), .A2(new_n334), .B1(new_n333), .B2(new_n257), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(KEYINPUT9), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n326), .A2(G200), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n328), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT10), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n336), .B1(new_n327), .B2(G169), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT67), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(KEYINPUT67), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(G179), .C2(new_n326), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n260), .ZN(new_n348));
  INV_X1    g0148(.A(new_n330), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n262), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n256), .A2(G1), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G20), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n348), .A2(new_n350), .B1(new_n352), .B2(new_n349), .ZN(new_n353));
  INV_X1    g0153(.A(new_n251), .ZN(new_n354));
  XNOR2_X1  g0154(.A(G58), .B(G68), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G20), .B1(G159), .B2(new_n243), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n213), .B2(new_n316), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT71), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT71), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n358), .C1(new_n213), .C2(new_n316), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n364), .B2(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n354), .B1(new_n365), .B2(KEYINPUT16), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT73), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n289), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n288), .A2(KEYINPUT73), .A3(G33), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n288), .B2(G33), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n286), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n213), .A2(new_n358), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n290), .A2(new_n209), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n373), .A2(new_n374), .B1(new_n375), .B2(new_n358), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n356), .B1(new_n376), .B2(new_n244), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n353), .B1(new_n366), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n323), .B1(G232), .B2(new_n324), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  OR2_X1    g0182(.A1(G223), .A2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G226), .B2(new_n318), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n382), .B1(new_n384), .B2(new_n290), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n283), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n381), .A2(G179), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n381), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT18), .B1(new_n380), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n290), .B2(new_n246), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n363), .B1(new_n392), .B2(new_n361), .ZN(new_n393));
  INV_X1    g0193(.A(new_n362), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n379), .A3(new_n251), .ZN(new_n397));
  INV_X1    g0197(.A(new_n353), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n390), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n311), .B1(new_n381), .B2(new_n386), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n381), .A2(new_n386), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(G190), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n404), .A4(new_n398), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n391), .A2(new_n401), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n260), .A2(G77), .A3(new_n262), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n257), .A2(new_n202), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n349), .A2(new_n243), .B1(new_n213), .B2(G77), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT15), .B(G87), .Z(new_n414));
  INV_X1    g0214(.A(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT68), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n413), .B1(new_n419), .B2(new_n247), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n412), .B1(new_n420), .B2(new_n251), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n316), .A2(G238), .A3(G1698), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n316), .A2(G232), .A3(new_n318), .ZN(new_n424));
  INV_X1    g0224(.A(G107), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(new_n316), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n283), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n323), .B1(G244), .B2(new_n324), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n422), .B1(G200), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n309), .B2(new_n429), .ZN(new_n431));
  AOI21_X1  g0231(.A(G169), .B1(new_n427), .B2(new_n428), .ZN(new_n432));
  OR3_X1    g0232(.A1(new_n421), .A2(new_n432), .A3(KEYINPUT69), .ZN(new_n433));
  INV_X1    g0233(.A(G179), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n427), .A2(new_n434), .A3(new_n428), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT69), .B1(new_n421), .B2(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n315), .A2(new_n347), .A3(new_n409), .A4(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(G1698), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(new_n318), .ZN(new_n441));
  INV_X1    g0241(.A(G294), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n440), .B(new_n441), .C1(new_n286), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n283), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G41), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n454));
  OAI211_X1 g0254(.A(G264), .B(new_n273), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n454), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(new_n450), .A3(new_n452), .A4(new_n269), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n444), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n388), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G179), .B2(new_n458), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n246), .A2(KEYINPUT23), .A3(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G116), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT84), .B1(new_n462), .B2(G20), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT84), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n209), .A3(G33), .A4(G116), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(G20), .B2(new_n425), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n461), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n246), .A2(new_n316), .A3(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT22), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT22), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n246), .A2(new_n316), .A3(new_n472), .A4(G87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n251), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n286), .A2(G1), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n257), .A2(new_n251), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n425), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT25), .B1(new_n257), .B2(new_n425), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n483), .A2(new_n425), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n460), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n354), .B1(new_n476), .B2(new_n478), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n458), .A2(G200), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n444), .A2(new_n455), .A3(G190), .A4(new_n457), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n490), .A2(new_n493), .A3(new_n487), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT85), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n493), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n480), .A2(new_n496), .A3(new_n488), .ZN(new_n497));
  INV_X1    g0297(.A(new_n458), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n434), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(new_n459), .C1(new_n490), .C2(new_n487), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n249), .A2(new_n250), .B1(G20), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n286), .A2(G97), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n505), .B1(new_n213), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n505), .B(KEYINPUT20), .C1(new_n213), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n352), .A2(G116), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n482), .B2(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(G270), .B(new_n273), .C1(new_n453), .C2(new_n454), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n316), .A2(G264), .A3(G1698), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n316), .A2(G257), .A3(new_n318), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n290), .A2(G303), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n434), .B1(new_n521), .B2(new_n283), .ZN(new_n522));
  AND4_X1   g0322(.A1(new_n457), .A2(new_n516), .A3(new_n517), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n283), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(new_n457), .A3(new_n517), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G169), .A3(new_n516), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT21), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n516), .A3(new_n528), .A4(G169), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n523), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n516), .B1(new_n525), .B2(G200), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n309), .B2(new_n525), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n439), .A2(new_n503), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT78), .A2(G250), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n446), .A2(new_n267), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G250), .ZN(new_n538));
  OAI22_X1  g0338(.A1(KEYINPUT78), .A2(new_n538), .B1(new_n445), .B2(G1), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n273), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n462), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G238), .A2(G1698), .ZN(new_n542));
  INV_X1    g0342(.A(G244), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(G1698), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n544), .B2(new_n316), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n540), .B1(new_n545), .B2(new_n282), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT79), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(KEYINPUT79), .B(new_n540), .C1(new_n545), .C2(new_n282), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(G190), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT81), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n548), .A2(new_n552), .A3(G190), .A4(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n210), .A2(new_n212), .A3(G33), .A4(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT80), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(KEYINPUT19), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(KEYINPUT80), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n246), .A2(new_n316), .A3(G68), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g0365(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n293), .B1(new_n559), .B2(new_n561), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n246), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n251), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n419), .A2(new_n257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n482), .A2(G87), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n548), .A2(new_n549), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(new_n311), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n551), .A2(KEYINPUT82), .A3(new_n553), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n556), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n373), .A2(new_n374), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n375), .A2(new_n358), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n425), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT6), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n581), .A2(new_n292), .A3(G107), .ZN(new_n582));
  XNOR2_X1  g0382(.A(G97), .B(G107), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n243), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n584), .A2(new_n246), .B1(new_n202), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n251), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n352), .A2(G97), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n482), .B2(G97), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n587), .A2(KEYINPUT74), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT74), .B1(new_n587), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT77), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n287), .A2(new_n289), .A3(G244), .A4(new_n318), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n507), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT75), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n596), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n282), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(new_n273), .C1(new_n453), .C2(new_n454), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n457), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n593), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n595), .A2(new_n596), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT75), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n595), .A2(new_n596), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n594), .A2(new_n507), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n600), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n283), .ZN(new_n611));
  INV_X1    g0411(.A(new_n603), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT77), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n604), .A2(G190), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n311), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n592), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n601), .A2(new_n593), .A3(new_n603), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT77), .B1(new_n611), .B2(new_n612), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n388), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n612), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(G179), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n587), .A2(new_n589), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n573), .A2(G169), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n548), .A2(new_n434), .A3(new_n549), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n482), .A2(new_n416), .A3(new_n418), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n569), .A2(new_n628), .A3(new_n570), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n577), .A2(new_n617), .A3(new_n625), .A4(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT83), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n604), .A2(new_n613), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n622), .B1(new_n636), .B2(new_n388), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n590), .A2(new_n591), .A3(new_n615), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n637), .A2(new_n624), .B1(new_n638), .B2(new_n614), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n574), .B1(new_n554), .B2(new_n555), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n631), .B1(new_n640), .B2(new_n576), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(KEYINPUT83), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n535), .B1(new_n635), .B2(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n307), .A2(new_n437), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n407), .A2(new_n408), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n314), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n399), .B(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n342), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n346), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(G169), .B1(new_n604), .B2(new_n613), .ZN(new_n652));
  INV_X1    g0452(.A(new_n624), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n652), .A2(new_n622), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n577), .A2(new_n654), .A3(new_n632), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n546), .A2(new_n388), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n627), .A2(new_n629), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n546), .A2(G200), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n551), .B2(new_n553), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n494), .A2(new_n662), .A3(new_n658), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n500), .A2(new_n530), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n625), .A3(new_n617), .A4(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n661), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n658), .B1(new_n554), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n590), .A2(new_n591), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(new_n637), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n656), .A2(new_n659), .A3(new_n665), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n439), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n651), .A2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n246), .A2(new_n674), .A3(new_n351), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n246), .A2(new_n351), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(G213), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n516), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n534), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n530), .B2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n684), .B1(new_n490), .B2(new_n487), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n503), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n684), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n500), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n489), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n684), .A2(new_n530), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n503), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(G399));
  NAND2_X1  g0499(.A1(new_n206), .A2(new_n451), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n261), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n566), .A2(new_n504), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n216), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n702), .A2(new_n704), .B1(new_n705), .B2(new_n701), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT28), .Z(new_n707));
  NAND4_X1  g0507(.A1(new_n495), .A2(new_n534), .A3(new_n502), .A4(new_n693), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n633), .A2(new_n634), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT83), .B1(new_n639), .B2(new_n641), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n573), .A2(new_n498), .A3(new_n517), .A4(new_n522), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n636), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n548), .A2(new_n522), .A3(new_n549), .A4(new_n517), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n458), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n604), .A4(new_n613), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n546), .A2(new_n434), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n621), .A2(new_n458), .A3(new_n525), .A4(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n684), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n689), .B1(new_n712), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT88), .ZN(new_n728));
  AND4_X1   g0528(.A1(new_n669), .A2(new_n667), .A3(new_n637), .A4(new_n668), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(KEYINPUT26), .B2(new_n655), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n664), .A2(new_n497), .A3(new_n667), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n658), .B1(new_n731), .B2(new_n639), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n684), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n728), .B1(new_n733), .B2(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n671), .A2(new_n693), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(KEYINPUT88), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n667), .A2(new_n637), .A3(new_n668), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT26), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n655), .B2(KEYINPUT26), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n664), .A2(new_n497), .A3(new_n667), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n617), .A2(new_n625), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n659), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT29), .B(new_n693), .C1(new_n741), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n727), .B1(new_n738), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n707), .B1(new_n746), .B2(G1), .ZN(G364));
  XOR2_X1   g0547(.A(new_n690), .B(KEYINPUT89), .Z(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n213), .A2(new_n256), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G45), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n702), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n752), .C1(G330), .C2(new_n687), .ZN(new_n753));
  INV_X1    g0553(.A(new_n752), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n316), .A2(new_n206), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n206), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n241), .A2(G45), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n290), .A2(new_n206), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n445), .B2(new_n705), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n250), .B1(G20), .B2(new_n388), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT90), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n754), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n434), .A2(new_n311), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT93), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(new_n246), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n246), .A2(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n434), .A2(new_n309), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n213), .A2(G200), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n775), .A2(G294), .B1(G326), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n773), .A2(new_n434), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT96), .Z(new_n784));
  NAND2_X1  g0584(.A1(new_n770), .A2(new_n772), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n311), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n772), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n786), .A2(G329), .B1(new_n789), .B2(G283), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(G20), .A3(G190), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n790), .B(new_n290), .C1(new_n791), .C2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n773), .A2(new_n434), .A3(new_n311), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G322), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n213), .A2(new_n311), .A3(new_n776), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT91), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n799), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n805), .A2(G58), .B1(new_n781), .B2(G77), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n785), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n797), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n244), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n812), .A2(new_n813), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n774), .A2(new_n292), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n795), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n290), .B1(new_n820), .B2(G87), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n789), .A2(G107), .B1(G50), .B2(new_n778), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n810), .A2(new_n819), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n784), .A2(new_n807), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n768), .B1(new_n825), .B2(new_n765), .ZN(new_n826));
  INV_X1    g0626(.A(new_n764), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n687), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n753), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND4_X1  g0630(.A1(new_n680), .A2(G343), .A3(new_n422), .A4(new_n681), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n431), .A2(new_n437), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n436), .A2(new_n435), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n684), .A2(new_n833), .A3(new_n422), .A4(new_n433), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n733), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n671), .A2(new_n693), .A3(new_n835), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT98), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n838), .ZN(new_n841));
  INV_X1    g0641(.A(new_n727), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT99), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n841), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n727), .B1(new_n844), .B2(new_n839), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n843), .A2(new_n752), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n844), .A2(new_n839), .A3(new_n727), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT99), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n832), .A2(new_n834), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n762), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n765), .A2(new_n762), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n754), .B1(G77), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n290), .B1(new_n777), .B2(new_n791), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n854), .B(new_n818), .C1(G116), .C2(new_n781), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n789), .A2(G87), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n856), .B1(new_n780), .B2(new_n785), .C1(new_n425), .C2(new_n795), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G294), .B2(new_n805), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n797), .A2(KEYINPUT97), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n797), .A2(KEYINPUT97), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n855), .B(new_n858), .C1(new_n859), .C2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n781), .A2(G159), .B1(G137), .B2(new_n778), .ZN(new_n864));
  INV_X1    g0664(.A(G150), .ZN(new_n865));
  INV_X1    g0665(.A(G143), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n865), .B2(new_n815), .C1(new_n866), .C2(new_n806), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT34), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n786), .A2(G132), .B1(new_n789), .B2(G68), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(new_n316), .C1(new_n333), .C2(new_n795), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G58), .B2(new_n775), .ZN(new_n872));
  INV_X1    g0672(.A(new_n867), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(KEYINPUT34), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n863), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n853), .B1(new_n875), .B2(new_n765), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n846), .A2(new_n848), .B1(new_n850), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(G384));
  INV_X1    g0678(.A(G58), .ZN(new_n879));
  OAI21_X1  g0679(.A(G77), .B1(new_n879), .B2(new_n244), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n880), .A2(new_n216), .B1(G50), .B2(new_n244), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n256), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT100), .Z(new_n883));
  NOR2_X1   g0683(.A1(new_n292), .A2(new_n425), .ZN(new_n884));
  NOR2_X1   g0684(.A1(G97), .A2(G107), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n581), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n582), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n504), .B(new_n215), .C1(new_n888), .C2(KEYINPUT35), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(KEYINPUT35), .B2(new_n888), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT36), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n395), .A2(new_n356), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n378), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n353), .B1(new_n366), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n405), .B1(new_n896), .B2(new_n682), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n390), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n399), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n680), .A2(new_n681), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n397), .A2(new_n398), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n900), .A2(new_n903), .A3(new_n904), .A4(new_n405), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n896), .A2(new_n682), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n409), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT38), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT38), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n900), .A2(new_n903), .A3(new_n405), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  INV_X1    g0715(.A(new_n903), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n915), .A2(new_n905), .B1(new_n409), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n912), .B(new_n913), .C1(KEYINPUT38), .C2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n911), .A2(KEYINPUT101), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n306), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n303), .A3(new_n300), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n264), .A3(new_n693), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n899), .A2(new_n905), .ZN(new_n925));
  INV_X1    g0725(.A(new_n907), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n647), .B2(new_n645), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n912), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT101), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT39), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n919), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n647), .A2(new_n901), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n684), .A2(new_n264), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n307), .A2(new_n314), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n307), .B2(new_n314), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n437), .A2(new_n684), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n837), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n933), .B1(new_n939), .B2(new_n929), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n745), .A2(new_n439), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n650), .B1(new_n738), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n941), .B(new_n943), .Z(new_n944));
  OAI21_X1  g0744(.A(new_n835), .B1(new_n935), .B2(new_n936), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n712), .B2(new_n726), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n929), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n399), .B1(new_n380), .B2(new_n404), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n904), .B1(new_n949), .B2(new_n903), .ZN(new_n950));
  INV_X1    g0750(.A(new_n905), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n903), .B1(new_n647), .B2(new_n645), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n924), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n948), .B1(new_n954), .B2(new_n912), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n947), .A2(new_n948), .B1(new_n955), .B2(new_n946), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n712), .A2(new_n726), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(new_n439), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n689), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n958), .B2(new_n956), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n944), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n261), .B2(new_n750), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n944), .A2(new_n960), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n893), .B1(new_n962), .B2(new_n963), .ZN(G367));
  INV_X1    g0764(.A(new_n572), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n684), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT102), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n658), .B2(new_n662), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n658), .B2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT103), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n684), .A2(new_n668), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(new_n637), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n743), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n698), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT42), .ZN(new_n978));
  INV_X1    g0778(.A(new_n976), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n654), .B1(new_n979), .B2(new_n489), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT104), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n693), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n980), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n972), .A2(KEYINPUT105), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n971), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n987), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT105), .B1(new_n972), .B2(new_n985), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n695), .A2(new_n976), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n991), .B(new_n992), .Z(new_n993));
  NAND2_X1  g0793(.A1(new_n751), .A2(G1), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n698), .A2(new_n696), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n976), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n976), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n695), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n698), .B1(new_n694), .B2(new_n697), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1004), .A2(new_n689), .A3(new_n688), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n749), .B2(new_n1004), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n746), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n746), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n700), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n995), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n993), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n316), .B1(new_n777), .B2(new_n866), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n774), .A2(new_n244), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G50), .C2(new_n781), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n786), .A2(G137), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n789), .A2(G77), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n879), .C2(new_n795), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G150), .B2(new_n805), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1017), .B(new_n1021), .C1(new_n811), .C2(new_n862), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n820), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT108), .Z(new_n1024));
  OAI22_X1  g0824(.A1(new_n859), .A2(new_n782), .B1(new_n774), .B2(new_n425), .ZN(new_n1025));
  INV_X1    g0825(.A(G317), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n290), .B1(new_n785), .B2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n788), .A2(new_n292), .B1(new_n780), .B2(new_n777), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1024), .B(new_n1029), .C1(new_n442), .C2(new_n862), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT46), .B1(new_n820), .B2(G116), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT109), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT109), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n791), .C2(new_n806), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1022), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT110), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT47), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n765), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n766), .B1(new_n419), .B2(new_n206), .C1(new_n233), .C2(new_n759), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n754), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n764), .B2(new_n971), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1014), .A2(new_n1042), .ZN(G387));
  OR2_X1    g0843(.A1(new_n694), .A2(new_n827), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n704), .A2(new_n755), .B1(G107), .B2(new_n206), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n759), .B1(new_n230), .B2(G45), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n445), .B1(new_n244), .B2(new_n202), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n703), .B2(KEYINPUT111), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n349), .A2(KEYINPUT50), .A3(new_n333), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT50), .B1(new_n349), .B2(new_n333), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1048), .B1(KEYINPUT111), .B2(new_n703), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1045), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n754), .B1(new_n1052), .B2(new_n767), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n774), .A2(new_n419), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n290), .B(new_n1054), .C1(G97), .C2(new_n789), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G68), .A2(new_n781), .B1(new_n797), .B2(new_n349), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n805), .A2(G50), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n795), .A2(new_n202), .B1(new_n811), .B2(new_n777), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G150), .B2(new_n786), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n316), .B1(new_n786), .B2(G326), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n774), .A2(new_n859), .B1(new_n442), .B2(new_n795), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n781), .A2(G303), .B1(G322), .B2(new_n778), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n1026), .B2(new_n806), .C1(new_n862), .C2(new_n780), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1061), .B1(new_n504), .B2(new_n788), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1060), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1053), .B1(new_n1071), .B2(new_n765), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1006), .A2(new_n994), .B1(new_n1044), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1007), .A2(new_n701), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1006), .A2(new_n746), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(G393));
  NAND2_X1  g0876(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1008), .A2(new_n701), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1003), .A2(new_n995), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n976), .A2(new_n764), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n238), .A2(new_n206), .A3(new_n290), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n766), .B1(new_n292), .B2(new_n206), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n754), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n805), .A2(G311), .B1(G317), .B2(new_n778), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n442), .A2(new_n782), .B1(new_n774), .B2(new_n504), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n290), .B1(new_n788), .B2(new_n425), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n795), .A2(new_n859), .B1(new_n785), .B2(new_n800), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1085), .B(new_n1089), .C1(new_n791), .C2(new_n862), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n775), .A2(G77), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n330), .B2(new_n782), .C1(new_n862), .C2(new_n333), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT112), .Z(new_n1093));
  AOI22_X1  g0893(.A1(new_n805), .A2(G159), .B1(G150), .B2(new_n778), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  AOI22_X1  g0895(.A1(new_n820), .A2(G68), .B1(new_n786), .B2(G143), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1095), .A2(new_n316), .A3(new_n856), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1090), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1083), .B1(new_n1098), .B2(new_n765), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1078), .A2(new_n1100), .A3(KEYINPUT113), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT113), .B1(new_n1078), .B2(new_n1100), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(new_n937), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n727), .A2(new_n835), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT114), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n837), .A2(new_n938), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1106), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n919), .A2(new_n931), .B1(new_n1112), .B2(new_n922), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n693), .B(new_n835), .C1(new_n741), .C2(new_n744), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n937), .B1(new_n1114), .B2(new_n938), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n912), .B1(new_n917), .B2(KEYINPUT38), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n922), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1107), .A2(new_n1108), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n708), .B1(new_n635), .B2(new_n642), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n724), .A2(new_n725), .ZN(new_n1121));
  OAI211_X1 g0921(.A(G330), .B(new_n835), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n937), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1114), .A2(new_n938), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1106), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n923), .B1(new_n954), .B2(new_n912), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1123), .A2(KEYINPUT114), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(KEYINPUT101), .B(new_n913), .C1(new_n928), .C2(new_n912), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n930), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n918), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n939), .A2(new_n923), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1109), .B(new_n1127), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1119), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT88), .B1(new_n735), .B2(new_n736), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n728), .B(KEYINPUT29), .C1(new_n671), .C2(new_n693), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n942), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n727), .A2(new_n439), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n651), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT115), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1136), .A2(KEYINPUT115), .A3(new_n651), .A4(new_n1137), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1106), .B1(new_n727), .B2(new_n835), .ZN(new_n1142));
  OAI211_X1 g0942(.A(KEYINPUT116), .B(new_n1111), .C1(new_n1142), .C2(new_n1123), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1122), .A2(new_n937), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1107), .A2(new_n938), .A3(new_n1144), .A4(new_n1114), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1107), .A2(new_n1144), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT116), .B1(new_n1147), .B2(new_n1111), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1140), .B(new_n1141), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n700), .B1(new_n1133), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1133), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1130), .A2(new_n763), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n786), .A2(G125), .B1(G128), .B2(new_n778), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n316), .C1(new_n333), .C2(new_n788), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n775), .A2(G159), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT53), .B1(new_n795), .B2(new_n865), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n820), .A2(G150), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1157), .B1(KEYINPUT53), .B2(new_n1158), .C1(new_n782), .C2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1154), .B(new_n1160), .C1(G132), .C2(new_n805), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n862), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(G137), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(G107), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n789), .A2(G68), .B1(G283), .B2(new_n778), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n442), .B2(new_n785), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n316), .B1(new_n820), .B2(G87), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1091), .B(new_n1167), .C1(new_n292), .C2(new_n782), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(G116), .C2(new_n805), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1161), .A2(new_n1163), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n765), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n754), .B1(new_n349), .B2(new_n852), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1152), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1119), .A2(new_n1132), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n994), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1151), .A2(new_n1175), .ZN(G378));
  AOI21_X1  g0976(.A(KEYINPUT115), .B1(new_n943), .B2(new_n1137), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1141), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1133), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1147), .A2(new_n1111), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT116), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1183), .B1(new_n1174), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1182), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n909), .A2(new_n910), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n307), .A2(new_n314), .A3(new_n934), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n264), .B(new_n684), .C1(new_n921), .C2(new_n313), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n849), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n948), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n946), .A2(KEYINPUT40), .A3(new_n1116), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(G330), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n901), .A2(new_n336), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n347), .B(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1197), .A2(new_n1198), .A3(G330), .A4(new_n1203), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n932), .A3(new_n940), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT119), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1203), .B1(new_n956), .B2(G330), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1206), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n941), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT120), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT120), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n941), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1209), .A2(new_n1213), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n941), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1215), .B1(new_n1214), .B2(new_n941), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1212), .A2(new_n1207), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT57), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1226));
  AOI211_X1 g1026(.A(KEYINPUT121), .B(new_n1183), .C1(new_n1174), .C2(new_n1187), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n701), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1223), .A2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n789), .A2(G58), .B1(G116), .B2(new_n778), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n859), .B2(new_n785), .C1(new_n806), .C2(new_n425), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n419), .A2(new_n782), .B1(new_n815), .B2(new_n292), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n316), .A2(G41), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n795), .B2(new_n202), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1016), .A4(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT58), .Z(new_n1237));
  OAI21_X1  g1037(.A(new_n333), .B1(G33), .B2(G41), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n778), .A2(G125), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n795), .A2(new_n1159), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(G132), .C2(new_n797), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n775), .A2(G150), .B1(G137), .B2(new_n781), .ZN(new_n1242));
  INV_X1    g1042(.A(G128), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1242), .C1(new_n1243), .C2(new_n806), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT117), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n286), .B(new_n451), .C1(new_n788), .C2(new_n811), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G124), .B2(new_n786), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT59), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1237), .B1(new_n1234), .B2(new_n1238), .C1(new_n1247), .C2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1171), .B1(new_n1252), .B2(KEYINPUT118), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(KEYINPUT118), .B2(new_n1252), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1254), .B(new_n754), .C1(G50), .C2(new_n852), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n762), .B2(new_n1204), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1222), .B2(new_n994), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1257), .ZN(G375));
  NAND2_X1  g1058(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1012), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1149), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n820), .A2(G97), .B1(new_n786), .B2(G303), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n442), .B2(new_n777), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G283), .B2(new_n805), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1019), .A2(new_n290), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1265), .B(new_n1054), .C1(G107), .C2(new_n781), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(new_n504), .C2(new_n862), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n316), .B1(new_n879), .B2(new_n788), .C1(new_n782), .C2(new_n865), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G50), .B2(new_n775), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n778), .A2(G132), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1270), .B1(new_n785), .B2(new_n1243), .C1(new_n795), .C2(new_n811), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G137), .B2(new_n805), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1269), .B(new_n1272), .C1(new_n862), .C2(new_n1159), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1171), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n752), .B(new_n1274), .C1(new_n244), .C2(new_n851), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n937), .A2(new_n762), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1180), .B2(new_n995), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1261), .A2(new_n1279), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT122), .Z(G381));
  NOR4_X1   g1081(.A1(G387), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1282));
  INV_X1    g1082(.A(G378), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1104), .A3(new_n1283), .ZN(new_n1284));
  OR3_X1    g1084(.A1(new_n1284), .A2(G375), .A3(G381), .ZN(G407));
  NAND2_X1  g1085(.A1(new_n683), .A2(G213), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT123), .Z(new_n1287));
  NAND4_X1  g1087(.A1(new_n1230), .A2(new_n1283), .A3(new_n1257), .A4(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(KEYINPUT124), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G407), .A2(new_n1289), .A3(G213), .ZN(G409));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G378), .B(new_n1257), .C1(new_n1223), .C2(new_n1229), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1256), .B1(new_n1224), .B2(new_n994), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1217), .B(new_n1221), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1012), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1283), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1287), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1180), .A2(new_n1183), .A3(KEYINPUT60), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1299), .A2(new_n701), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1259), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G384), .B1(new_n1303), .B2(new_n1279), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n877), .B(new_n1278), .C1(new_n1300), .C2(new_n1302), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT125), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1179), .B2(new_n1187), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1179), .A2(new_n1187), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1299), .A2(new_n701), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1279), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n877), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1303), .A2(G384), .A3(new_n1279), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1287), .A2(G2897), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1306), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1317), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1314), .A3(new_n1320), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1297), .A2(new_n1298), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1291), .B1(new_n1322), .B2(KEYINPUT61), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1287), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT126), .B(new_n1324), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1319), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1319), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(KEYINPUT62), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1323), .A2(new_n1327), .A3(new_n1329), .A4(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(G387), .A2(new_n1104), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(G390), .A2(new_n1014), .A3(new_n1042), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(G393), .B(new_n829), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1333), .A2(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1322), .A2(KEYINPUT61), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1330), .A2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1339), .A2(new_n1342), .A3(new_n1343), .A4(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1341), .A2(new_n1346), .ZN(G405));
  INV_X1    g1147(.A(new_n1319), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G375), .A2(new_n1283), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1349), .B2(new_n1292), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1349), .A2(new_n1292), .A3(new_n1348), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1340), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1350), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1339), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(G402));
endmodule


