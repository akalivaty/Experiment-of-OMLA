//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n461), .B1(new_n450), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n472), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n465), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n466), .A2(new_n467), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(new_n465), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n480), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(G124), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT72), .Z(G162));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n478), .B2(new_n479), .ZN(new_n494));
  AND2_X1   g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n465), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n478), .B2(new_n479), .ZN(new_n498));
  AND2_X1   g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n496), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(new_n509), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT73), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT74), .B(G88), .Z(new_n518));
  AOI21_X1  g093(.A(new_n507), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n520), .B2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n508), .A2(new_n509), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n510), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(KEYINPUT75), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(KEYINPUT75), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n517), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n520), .A2(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n511), .A2(new_n516), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(G90), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n538), .B1(new_n510), .B2(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT77), .ZN(G171));
  NAND2_X1  g118(.A1(new_n517), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT5), .B(G543), .Z(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n520), .A2(G43), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(G65), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(G65), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n522), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n510), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n516), .A2(new_n519), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n516), .A2(new_n566), .A3(G53), .A4(new_n519), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n562), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n540), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT78), .A4(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n568), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n517), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n520), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n522), .A2(G61), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(G73), .B2(G543), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n522), .A2(KEYINPUT80), .A3(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n510), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(G86), .A2(new_n517), .B1(new_n520), .B2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(G85), .A2(new_n517), .B1(new_n520), .B2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n590), .A2(KEYINPUT82), .A3(new_n510), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT82), .B1(new_n590), .B2(new_n510), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(G290));
  NAND3_X1  g168(.A1(new_n511), .A2(new_n516), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n546), .A2(new_n597), .B1(new_n598), .B2(new_n507), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI221_X1 g176(.A(KEYINPUT84), .B1(new_n598), .B2(new_n507), .C1(new_n546), .C2(new_n597), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(G651), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n563), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(new_n563), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n596), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G171), .B2(G868), .ZN(G284));
  XNOR2_X1  g185(.A(G284), .B(KEYINPUT85), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  AND3_X1   g190(.A1(new_n596), .A2(new_n603), .A3(new_n607), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n551), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n612), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n608), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n480), .A2(new_n473), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n490), .A2(G123), .ZN(new_n630));
  INV_X1    g205(.A(new_n481), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT88), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n632), .A2(KEYINPUT88), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n631), .A2(G135), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n627), .A2(G2100), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n629), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT89), .Z(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n652), .B2(new_n653), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  INV_X1    g238(.A(new_n660), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n658), .B(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n667), .B2(new_n664), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n664), .A3(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n674), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G160), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT24), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n692), .A2(G34), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n691), .B1(new_n692), .B2(G34), .ZN(new_n694));
  OAI22_X1  g269(.A1(new_n690), .A2(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G2084), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G5), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G171), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G1961), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT26), .Z(new_n703));
  NAND3_X1  g278(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G141), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n703), .B(new_n706), .C1(new_n707), .C2(new_n481), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G129), .B2(new_n490), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G32), .B(new_n712), .S(G29), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  AOI211_X1 g289(.A(new_n697), .B(new_n701), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT98), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT98), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G1961), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n698), .A2(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n551), .B2(new_n698), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1341), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n698), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n698), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT97), .B(G1966), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n718), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(G29), .A2(G33), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n631), .A2(G139), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n465), .C2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n691), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n691), .A2(G26), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  INV_X1    g314(.A(G140), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n465), .A2(G116), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n481), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G128), .B2(new_n490), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n739), .B1(new_n744), .B2(new_n691), .ZN(new_n745));
  INV_X1    g320(.A(G2067), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT30), .B(G28), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n748), .A2(new_n691), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n637), .B2(new_n691), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n695), .A2(new_n696), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n735), .C2(new_n734), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n737), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G27), .A2(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G164), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT99), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n698), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n726), .A2(new_n755), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n716), .A2(new_n717), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G29), .A2(G35), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G162), .B2(G29), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n616), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G4), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(G1348), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n776), .B(new_n777), .C1(new_n713), .C2(new_n714), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n771), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n698), .A2(G24), .ZN(new_n781));
  INV_X1    g356(.A(G290), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n698), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(G1986), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n691), .A2(G25), .ZN(new_n785));
  NOR2_X1   g360(.A1(G95), .A2(G2105), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT91), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n788));
  INV_X1    g363(.A(G131), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n787), .A2(new_n788), .B1(new_n481), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G119), .B2(new_n490), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(new_n691), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n783), .A2(G1986), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n698), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n698), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT33), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1976), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n698), .A2(G6), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G305), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n698), .A2(G22), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT92), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G303), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1971), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n801), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n784), .B(new_n796), .C1(new_n810), .C2(KEYINPUT34), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT36), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n780), .B1(new_n814), .B2(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n816), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n818), .A2(new_n779), .A3(new_n766), .ZN(G150));
  INV_X1    g394(.A(G860), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(new_n510), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n511), .A2(new_n516), .A3(G93), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n516), .A2(G55), .A3(new_n519), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n825), .B1(new_n824), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(new_n823), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n619), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n829), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n831), .A3(new_n551), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n616), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n821), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT102), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT102), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n820), .B1(new_n821), .B2(new_n839), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n829), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(G162), .B(G160), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT103), .ZN(new_n848));
  INV_X1    g423(.A(new_n637), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n847), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n637), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n712), .B(new_n504), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(new_n626), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n626), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n631), .A2(G142), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n465), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(G130), .B2(new_n490), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n791), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n744), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n856), .A2(new_n857), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n856), .B2(new_n857), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n854), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n871), .A2(new_n850), .A3(new_n853), .A4(new_n867), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(new_n836), .B(new_n621), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n877));
  NAND2_X1  g452(.A1(G299), .A2(KEYINPUT105), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n568), .A2(new_n879), .A3(new_n573), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n616), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n608), .A2(KEYINPUT105), .A3(G299), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n877), .B1(new_n883), .B2(KEYINPUT41), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n887), .A3(new_n882), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n876), .B(new_n885), .C1(new_n889), .C2(KEYINPUT106), .ZN(new_n890));
  INV_X1    g465(.A(new_n883), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n876), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G305), .B(G303), .ZN(new_n897));
  XNOR2_X1  g472(.A(G290), .B(G288), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n894), .B2(new_n895), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n892), .A4(KEYINPUT42), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n896), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n896), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(G868), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n829), .A2(new_n612), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n906), .ZN(G331));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND3_X1  g484(.A1(G171), .A2(new_n835), .A3(new_n833), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G171), .B1(new_n833), .B2(new_n835), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n911), .A2(new_n912), .A3(G286), .ZN(new_n913));
  NAND2_X1  g488(.A1(G301), .A2(new_n836), .ZN(new_n914));
  AOI21_X1  g489(.A(G168), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT106), .B1(new_n886), .B2(new_n888), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n913), .A2(new_n915), .B1(new_n916), .B2(new_n884), .ZN(new_n917));
  OAI21_X1  g492(.A(G286), .B1(new_n911), .B2(new_n912), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(G168), .A3(new_n910), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n891), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n899), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n873), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n899), .B1(new_n917), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n909), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n920), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n889), .B1(new_n919), .B2(new_n918), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n900), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(KEYINPUT43), .A3(new_n921), .A4(new_n873), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT44), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n922), .B2(new_n923), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(new_n909), .A3(new_n921), .A4(new_n873), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(G397));
  XNOR2_X1  g511(.A(new_n744), .B(new_n746), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n712), .B2(G1996), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n504), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n470), .A2(new_n475), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n939), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT45), .B1(new_n504), .B2(new_n940), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(KEYINPUT109), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n938), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n954), .A2(KEYINPUT110), .A3(new_n712), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n954), .B2(new_n712), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n791), .B(new_n793), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(G1986), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT113), .B(G8), .Z(new_n963));
  AND3_X1   g538(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(new_n948), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n945), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n724), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n941), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n941), .A2(KEYINPUT50), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT116), .B(G2084), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n969), .A2(new_n945), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n963), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(G168), .A2(new_n963), .ZN(new_n974));
  OR3_X1    g549(.A1(new_n973), .A2(KEYINPUT51), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n967), .A2(new_n972), .ZN(new_n976));
  INV_X1    g551(.A(new_n963), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT51), .B1(new_n978), .B2(G168), .ZN(new_n979));
  INV_X1    g554(.A(G8), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n967), .B2(new_n972), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(new_n974), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT114), .B(G1981), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n586), .A2(new_n587), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n587), .B(KEYINPUT115), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n586), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT49), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n586), .B2(new_n986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n584), .A2(KEYINPUT81), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n584), .A2(KEYINPUT81), .ZN(new_n993));
  AND4_X1   g568(.A1(new_n992), .A2(new_n993), .A3(new_n587), .A4(new_n984), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n945), .A2(new_n504), .A3(new_n940), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n977), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G8), .B1(new_n525), .B2(new_n526), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT111), .B(G1971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n966), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n969), .A2(new_n770), .A3(new_n945), .A4(new_n970), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n980), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n941), .A2(new_n968), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n504), .A2(new_n1009), .A3(new_n940), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n945), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2090), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n966), .B2(new_n1003), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1001), .B1(new_n1013), .B2(new_n963), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n798), .B2(G1976), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n997), .B1(G1976), .B2(new_n798), .ZN(new_n1017));
  MUX2_X1   g592(.A(new_n1015), .B(new_n1016), .S(new_n1017), .Z(new_n1018));
  NAND4_X1  g593(.A1(new_n999), .A2(new_n1007), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n983), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n966), .B2(G2078), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n969), .A2(new_n945), .A3(new_n970), .ZN(new_n1023));
  INV_X1    g598(.A(G1961), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1021), .A2(G2078), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n965), .A2(G40), .A3(G160), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT124), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1022), .A2(new_n1030), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(G171), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n965), .A2(new_n945), .A3(new_n1026), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1022), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(G301), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(G171), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n1033), .C1(G171), .C2(new_n1028), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1020), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT61), .ZN(new_n1042));
  NOR2_X1   g617(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT118), .Z(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(G299), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1048), .B(new_n1044), .C1(new_n568), .C2(new_n573), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT56), .B(G2072), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n965), .A2(KEYINPUT119), .A3(new_n945), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1011), .A2(new_n763), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n943), .A2(new_n945), .A3(new_n1056), .A4(new_n1053), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND4_X1   g634(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(new_n1057), .B1(new_n1011), .B2(new_n763), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1052), .B1(new_n1061), .B2(new_n1054), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1042), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n943), .A2(new_n953), .A3(new_n945), .A4(new_n1056), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  AND3_X1   g642(.A1(new_n996), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n996), .B2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1065), .B(KEYINPUT122), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1064), .B1(new_n1074), .B2(new_n551), .ZN(new_n1075));
  AOI211_X1 g650(.A(KEYINPUT59), .B(new_n619), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1063), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1061), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT61), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1061), .A2(new_n1080), .A3(new_n1054), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1054), .A2(new_n1059), .A3(new_n1055), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1052), .B1(new_n1082), .B2(KEYINPUT120), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1079), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT123), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1069), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n996), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT122), .B1(new_n1088), .B2(new_n1065), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1073), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n551), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1074), .A2(new_n1064), .A3(new_n551), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1082), .A2(KEYINPUT120), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1052), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1081), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1078), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1094), .A2(new_n1098), .A3(new_n1099), .A4(new_n1063), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n996), .A2(G2067), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1023), .B2(new_n775), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n608), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n608), .B1(new_n1102), .B2(KEYINPUT60), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1103), .A2(new_n1104), .B1(KEYINPUT60), .B2(new_n1102), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1085), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1097), .B1(new_n608), .B2(new_n1102), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1078), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1041), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n975), .B(KEYINPUT62), .C1(new_n979), .C2(new_n982), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT125), .ZN(new_n1111));
  OAI221_X1 g686(.A(KEYINPUT51), .B1(new_n981), .B2(new_n974), .C1(new_n978), .C2(G168), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT62), .A4(new_n975), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n983), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1019), .A2(new_n1038), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(G288), .A2(G1976), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n994), .B1(new_n999), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n999), .A2(new_n1018), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1120), .A2(new_n997), .B1(new_n1121), .B2(new_n1007), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1121), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n973), .A2(G168), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(new_n1007), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1019), .B2(new_n1125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1118), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n962), .B1(new_n1109), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n957), .A2(new_n959), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n950), .A2(G1986), .A3(G290), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT48), .Z(new_n1135));
  OAI21_X1  g710(.A(new_n952), .B1(new_n712), .B2(new_n937), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n954), .A2(KEYINPUT46), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n954), .A2(KEYINPUT46), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT47), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(KEYINPUT47), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1133), .A2(new_n1135), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n791), .A2(new_n793), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT126), .Z(new_n1145));
  AOI22_X1  g720(.A1(new_n957), .A2(new_n1145), .B1(new_n746), .B2(new_n744), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1146), .B2(new_n950), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1146), .A2(new_n1143), .A3(new_n950), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g726(.A1(new_n463), .A2(G227), .ZN(new_n1153));
  NOR3_X1   g727(.A1(G401), .A2(G229), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g728(.A1(new_n933), .A2(new_n1154), .A3(new_n874), .ZN(G225));
  INV_X1    g729(.A(G225), .ZN(G308));
endmodule


