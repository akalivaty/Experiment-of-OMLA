//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142,
    new_n1143, new_n1145;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g027(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n453));
  NAND3_X1  g028(.A1(new_n437), .A2(new_n438), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n456), .ZN(new_n460));
  INV_X1    g035(.A(new_n457), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n460), .A2(G2106), .B1(G567), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n467), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n470), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT68), .Z(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(new_n466), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n469), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(G124), .A2(new_n478), .B1(new_n479), .B2(G136), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n476), .A2(new_n480), .ZN(G162));
  NAND2_X1  g056(.A1(G114), .A2(G2104), .ZN(new_n482));
  INV_X1    g057(.A(G126), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n482), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n467), .A2(G138), .A3(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  INV_X1    g065(.A(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n469), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT70), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(G651), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n510), .A2(new_n506), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  NAND2_X1  g091(.A1(G63), .A2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n500), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n508), .A2(new_n500), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G89), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n508), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n505), .A2(KEYINPUT71), .A3(new_n507), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G51), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n514), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n520), .A2(new_n514), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n500), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  INV_X1    g108(.A(new_n519), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OR2_X1    g110(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n506), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n507), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n522), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n540), .A2(G543), .A3(new_n524), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n533), .B1(new_n534), .B2(new_n535), .C1(new_n541), .C2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(new_n541), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n500), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n506), .B1(new_n549), .B2(KEYINPUT73), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n550), .B1(KEYINPUT73), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n519), .A2(G81), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n546), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n540), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT74), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT74), .B1(new_n497), .B2(new_n499), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G78), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n521), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n523), .A2(KEYINPUT9), .A3(G53), .A4(new_n524), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n519), .A2(G91), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n562), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n538), .A2(new_n539), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n575), .A2(G91), .A3(new_n501), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n500), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(G65), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n567), .B2(new_n521), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n576), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n582), .A2(KEYINPUT75), .A3(new_n570), .A4(new_n562), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n574), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n545), .A2(G49), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT76), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n506), .B1(new_n500), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n519), .B2(G87), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n519), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n500), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n575), .A2(G48), .A3(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n519), .A2(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n599), .B1(new_n506), .B2(new_n600), .C1(new_n541), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n541), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n578), .A2(G66), .A3(new_n579), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n506), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n604), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G651), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n523), .A2(G54), .A3(new_n524), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n612), .A2(KEYINPUT77), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n534), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n610), .A2(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n603), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n603), .B1(new_n619), .B2(G868), .ZN(G321));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g197(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n619), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n479), .A2(G2104), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT13), .Z(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n479), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n478), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n469), .B2(G111), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n634), .A2(new_n635), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT79), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT81), .ZN(new_n647));
  INV_X1    g222(.A(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n650), .B2(new_n649), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n662), .A3(new_n658), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  INV_X1    g248(.A(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n670), .B1(new_n674), .B2(new_n668), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT83), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(KEYINPUT83), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n668), .B(KEYINPUT17), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n677), .C1(new_n674), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n670), .A3(new_n674), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n673), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n641), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2100), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT84), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  INV_X1    g272(.A(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n696), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT86), .B(G1986), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NOR2_X1   g280(.A1(G160), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  NOR2_X1   g282(.A1(KEYINPUT24), .A2(G34), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n706), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2084), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT99), .Z(new_n713));
  AND2_X1   g288(.A1(new_n705), .A2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n479), .A2(G141), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT95), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n478), .A2(G129), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n714), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT31), .B(G11), .Z(new_n728));
  INV_X1    g303(.A(G28), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT97), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n727), .B(new_n733), .C1(new_n705), .C2(new_n640), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n710), .A2(new_n711), .B1(new_n725), .B2(new_n726), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n479), .A2(G140), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n478), .A2(G128), .ZN(new_n737));
  NOR2_X1   g312(.A1(G104), .A2(G2105), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n705), .A2(G26), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2067), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n734), .A2(new_n735), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n554), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G1341), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(G1341), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n713), .A2(new_n746), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n747), .A2(G4), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n619), .B2(new_n747), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n752), .B1(G1348), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G21), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G168), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n755), .B(new_n759), .C1(G1348), .C2(new_n754), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT92), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n479), .A2(G139), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n764), .B(new_n765), .C1(new_n469), .C2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G33), .B(new_n767), .S(G29), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT93), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2072), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT94), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n705), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n705), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT100), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT29), .B(G2090), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n705), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n705), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n780), .C1(G2072), .C2(new_n769), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n747), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n747), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n760), .A2(new_n771), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n747), .A2(G23), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n587), .A2(new_n590), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n747), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G6), .A2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G305), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(new_n698), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n747), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n747), .ZN(new_n799));
  INV_X1    g374(.A(G1971), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n790), .A2(new_n791), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n792), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n478), .A2(G119), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT87), .Z(new_n807));
  OR2_X1    g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(G107), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n491), .B1(new_n809), .B2(G2105), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n479), .A2(G131), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n705), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G25), .B2(new_n705), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT88), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n815), .A2(new_n817), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n747), .A2(G24), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT89), .Z(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G290), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1986), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n804), .A2(new_n805), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n747), .A2(G20), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT23), .ZN(new_n831));
  INV_X1    g406(.A(G299), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n747), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G1956), .Z(new_n834));
  NAND4_X1  g409(.A1(new_n787), .A2(new_n828), .A3(new_n829), .A4(new_n834), .ZN(G150));
  INV_X1    g410(.A(G150), .ZN(G311));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n500), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G651), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n840), .B1(new_n534), .B2(new_n841), .C1(new_n541), .C2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n554), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n553), .A2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT38), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n619), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT101), .B(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n844), .A2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n494), .B(new_n740), .ZN(new_n858));
  INV_X1    g433(.A(new_n724), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n767), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n479), .A2(G142), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n478), .A2(G130), .ZN(new_n863));
  NOR2_X1   g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(new_n469), .B2(G118), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n812), .B(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(new_n632), .Z(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n861), .A2(new_n869), .ZN(new_n871));
  XNOR2_X1  g446(.A(G162), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT102), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n640), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n871), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(KEYINPUT103), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n878), .A2(new_n861), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n861), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n874), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n876), .B(new_n877), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g458(.A1(new_n789), .A2(G305), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G303), .ZN(new_n885));
  AOI21_X1  g460(.A(G305), .B1(new_n587), .B2(new_n590), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n885), .ZN(new_n889));
  NOR2_X1   g464(.A1(G288), .A2(new_n794), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n847), .B(new_n626), .Z(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(G299), .B2(new_n619), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(new_n619), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n617), .A2(new_n618), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n606), .A2(new_n609), .A3(new_n604), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT77), .B1(new_n612), .B2(new_n613), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n574), .A4(new_n583), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(G299), .B2(new_n619), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n896), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n906), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n896), .A2(new_n907), .A3(KEYINPUT105), .A4(new_n902), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n894), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n893), .A2(new_n905), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n893), .B1(new_n905), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n844), .A2(G868), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G295));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n917), .A2(new_n920), .A3(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G331));
  XOR2_X1   g498(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n924));
  INV_X1    g499(.A(new_n892), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n527), .A2(new_n528), .A3(G301), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G301), .B1(new_n527), .B2(new_n528), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n847), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n846), .A3(new_n845), .A4(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n908), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n911), .B2(KEYINPUT109), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n903), .A2(new_n936), .A3(new_n906), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n933), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n904), .A2(new_n932), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n925), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n913), .B2(new_n932), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n941), .B2(new_n892), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n909), .A2(new_n908), .B1(new_n903), .B2(new_n906), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n933), .B1(new_n945), .B2(new_n912), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n925), .B1(new_n946), .B2(new_n939), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n948), .B2(KEYINPUT108), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  AOI211_X1 g525(.A(new_n950), .B(new_n943), .C1(new_n942), .C2(new_n947), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n924), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n940), .A2(new_n942), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT44), .B(new_n953), .C1(new_n954), .C2(new_n943), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n494), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n488), .B2(new_n493), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G160), .A2(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n959), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(G1996), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n740), .B(G2067), .Z(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n859), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT126), .Z(new_n972));
  NOR2_X1   g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n724), .B(G1996), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n969), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n813), .A2(new_n816), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n976), .A2(new_n977), .B1(G2067), .B2(new_n740), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n965), .ZN(new_n979));
  OR3_X1    g554(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n813), .A2(new_n816), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n969), .A2(new_n982), .A3(new_n975), .A4(new_n977), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n980), .A2(new_n981), .B1(new_n966), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n980), .A2(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n974), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G40), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n470), .A2(new_n472), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n961), .A2(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n990), .A2(KEYINPUT111), .A3(G8), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n990), .B2(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(G305), .B(G1981), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT49), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n991), .B2(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n789), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n794), .A2(new_n698), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n991), .A2(new_n992), .B1(G288), .B2(new_n997), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT52), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n789), .B2(G1976), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1002), .B(new_n996), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n958), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n964), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n964), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n958), .A2(new_n960), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n800), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1007), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT55), .Z(new_n1020));
  AND2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1000), .B1(new_n1006), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(KEYINPUT113), .A2(KEYINPUT63), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n989), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n758), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1966), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1011), .A2(new_n711), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(G8), .A3(G168), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1024), .A2(new_n1006), .A3(new_n1025), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(KEYINPUT113), .A2(KEYINPUT63), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1005), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1025), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1022), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n1044));
  AOI211_X1 g619(.A(new_n1008), .B(G1384), .C1(new_n488), .C2(new_n493), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n989), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n1032), .A2(KEYINPUT112), .B1(new_n1046), .B2(G2084), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1048));
  OAI21_X1  g623(.A(G8), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G168), .A2(new_n1007), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(KEYINPUT51), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(G8), .C1(new_n1035), .C2(G286), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1035), .A2(new_n1055), .A3(new_n1050), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n1035), .B2(new_n1050), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1052), .B(new_n1054), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1014), .A2(new_n1015), .A3(new_n779), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1061), .A2(new_n1062), .B1(new_n1046), .B2(new_n785), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT56), .B(G2072), .Z(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT114), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1014), .A2(new_n1015), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1011), .B2(G1956), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n572), .B(KEYINPUT57), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n990), .A2(G2067), .ZN(new_n1074));
  INV_X1    g649(.A(G1348), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1046), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n901), .B2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT115), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1011), .A2(G1348), .B1(G2067), .B2(new_n990), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n619), .A2(new_n1081), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n619), .A2(KEYINPUT121), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1086), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n619), .A2(KEYINPUT121), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1073), .A2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1095), .B(KEYINPUT61), .C1(new_n1083), .C2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1078), .B(new_n1073), .C1(new_n1094), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n990), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT116), .B1(new_n1016), .B2(G1996), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1016), .A2(KEYINPUT116), .A3(G1996), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n554), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1109), .B2(KEYINPUT59), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1085), .B1(new_n1100), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT53), .B1(new_n1116), .B2(new_n779), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1116), .B2(new_n779), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1014), .B(new_n1118), .C1(new_n959), .C2(new_n963), .ZN(new_n1119));
  AOI21_X1  g694(.A(G301), .B1(new_n1063), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1120), .A2(KEYINPUT125), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1064), .A2(G171), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(KEYINPUT125), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1063), .A2(new_n1126), .A3(G301), .A4(new_n1119), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1065), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1063), .A2(G301), .A3(new_n1119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT124), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1124), .A2(KEYINPUT54), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1067), .B1(new_n1115), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1059), .B1(KEYINPUT62), .B2(new_n1066), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1041), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1043), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(G290), .B(new_n823), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n966), .B1(new_n983), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n987), .B1(new_n1136), .B2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g714(.A1(new_n949), .A2(new_n951), .ZN(new_n1141));
  NOR3_X1   g715(.A1(G229), .A2(new_n463), .A3(G227), .ZN(new_n1142));
  NAND3_X1  g716(.A1(new_n666), .A2(new_n882), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1143), .ZN(G308));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1145));
  OAI21_X1  g719(.A(new_n1145), .B1(new_n951), .B2(new_n949), .ZN(G225));
endmodule


