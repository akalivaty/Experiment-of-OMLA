//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n459), .B2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n460), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n459), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n461), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n466), .A2(new_n472), .A3(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n471), .A2(G136), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT66), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(G2105), .A3(new_n469), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n477), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(G162));
  NAND4_X1  g061(.A1(new_n468), .A2(G138), .A3(new_n465), .A4(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n460), .A2(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR4_X1   g068(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n493), .A4(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n497), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT70), .B1(new_n497), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n469), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n460), .B2(new_n467), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n503), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT72), .A3(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT73), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(new_n523), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n516), .A2(new_n520), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n518), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n521), .A2(new_n539), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n518), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n521), .A2(new_n545), .B1(new_n523), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT76), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n521), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n516), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT78), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n565), .A3(G651), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n558), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n523), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n569), .B2(new_n570), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n567), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n534), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n530), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT79), .ZN(G288));
  AOI22_X1  g159(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n585), .A2(KEYINPUT80), .A3(new_n518), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT80), .B1(new_n585), .B2(new_n518), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n534), .A2(G86), .B1(new_n530), .B2(G48), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G305));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n521), .A2(new_n590), .B1(new_n523), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n518), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n534), .A2(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n560), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT82), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  XOR2_X1   g188(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  INV_X1    g191(.A(new_n548), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n611), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n608), .A2(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n471), .A2(G135), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n465), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n479), .A2(G123), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n463), .A2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(G2100), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n632), .B2(new_n631), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n637), .ZN(G156));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT16), .B(G1341), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n644), .A2(new_n650), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(KEYINPUT17), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n662), .C1(new_n663), .C2(new_n659), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n662), .A2(KEYINPUT18), .A3(new_n658), .ZN(new_n665));
  OAI21_X1  g240(.A(KEYINPUT18), .B1(new_n662), .B2(new_n658), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT86), .B(G2096), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n673), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT87), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(KEYINPUT87), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1991), .ZN(new_n688));
  INV_X1    g263(.A(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT29), .Z(new_n701));
  INV_X1    g276(.A(G2090), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT97), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n698), .A2(G33), .ZN(new_n705));
  NAND2_X1  g280(.A1(G115), .A2(G2104), .ZN(new_n706));
  INV_X1    g281(.A(G127), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n492), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT94), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n473), .A2(G103), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  INV_X1    g287(.A(G139), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n470), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(KEYINPUT93), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(KEYINPUT93), .B2(new_n714), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n705), .B1(new_n716), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n719));
  INV_X1    g294(.A(G26), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G29), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G128), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n471), .A2(G140), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n465), .A2(G116), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n722), .B1(new_n727), .B2(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n721), .B1(new_n728), .B2(new_n719), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n718), .A2(G2072), .B1(G2067), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G2067), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(G4), .A2(G16), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n608), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n698), .B1(KEYINPUT24), .B2(G34), .ZN(new_n737));
  OAI22_X1  g312(.A1(G160), .A2(new_n698), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2084), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT30), .B(G28), .Z(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  AND2_X1   g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n739), .B1(G29), .B2(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G21), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G168), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1966), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n738), .A2(G2084), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n623), .A2(G29), .A3(new_n627), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(G171), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G5), .B2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n743), .A2(new_n746), .A3(new_n747), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n548), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(G19), .ZN(new_n758));
  INV_X1    g333(.A(G1341), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n758), .A2(new_n759), .B1(new_n751), .B2(new_n753), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n760), .B1(new_n759), .B2(new_n758), .C1(new_n749), .C2(new_n748), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G2072), .B2(new_n718), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n731), .A2(new_n735), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n756), .A2(G20), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n764), .B(new_n765), .C1(G299), .C2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT98), .B(G1956), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n698), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n698), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G2078), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G32), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n471), .A2(G141), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n479), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(G105), .B2(new_n473), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n774), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT95), .Z(new_n782));
  AOI21_X1  g357(.A(new_n773), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n771), .A2(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n763), .A2(new_n769), .A3(new_n772), .A4(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n704), .B(new_n788), .C1(new_n702), .C2(new_n701), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(new_n583), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n756), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n756), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G1971), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(G1971), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n756), .A2(G6), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G305), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n479), .A2(G119), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n471), .A2(G131), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n465), .A2(G107), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(G29), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT90), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n756), .A2(G24), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n597), .B2(new_n756), .ZN(new_n818));
  INV_X1    g393(.A(G1986), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n806), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT92), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n789), .A2(new_n825), .ZN(G311));
  XNOR2_X1  g401(.A(G311), .B(KEYINPUT99), .ZN(G150));
  NAND2_X1  g402(.A1(new_n608), .A2(G559), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n518), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n521), .A2(new_n833), .B1(new_n523), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n548), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n617), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n830), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XOR2_X1   g421(.A(G162), .B(G160), .Z(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n628), .Z(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  MUX2_X1   g424(.A(new_n782), .B(new_n781), .S(new_n716), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n509), .B(new_n727), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n479), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n471), .A2(G142), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n465), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n811), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT100), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n631), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n849), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n850), .B(new_n851), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n861), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n848), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT101), .B1(new_n864), .B2(new_n861), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n847), .B(new_n628), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n853), .A2(new_n862), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(G395));
  XNOR2_X1  g449(.A(new_n619), .B(new_n841), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n607), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n602), .A2(new_n606), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(new_n567), .A3(new_n575), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n881), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n597), .A2(new_n583), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n594), .A2(new_n583), .A3(new_n596), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G305), .B(G166), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G290), .A2(new_n791), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(KEYINPUT103), .A3(new_n889), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n891), .A3(new_n892), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT42), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n886), .A2(new_n898), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n611), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n836), .A2(G868), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT104), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  OR2_X1    g480(.A1(new_n901), .A2(new_n902), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  NAND2_X1  g482(.A1(G286), .A2(G171), .ZN(new_n908));
  NAND2_X1  g483(.A1(G168), .A2(G301), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n841), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n840), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n883), .A2(new_n884), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n910), .A3(new_n879), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT105), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n910), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n885), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n920), .A3(new_n897), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n913), .A2(new_n915), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n897), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n867), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n907), .B1(new_n924), .B2(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n867), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n897), .B1(new_n916), .B2(new_n920), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n925), .B1(KEYINPUT43), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n923), .A2(new_n931), .A3(new_n921), .A4(new_n867), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT106), .B1(new_n933), .B2(new_n907), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n935));
  AOI211_X1 g510(.A(new_n935), .B(KEYINPUT44), .C1(new_n930), .C2(new_n932), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n929), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n939), .B(new_n929), .C1(new_n934), .C2(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(G397));
  AND2_X1   g516(.A1(G160), .A2(G40), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n509), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(KEYINPUT110), .B(G1384), .C1(new_n496), .C2(new_n508), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G8), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G305), .A2(G1981), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n586), .A2(new_n694), .A3(new_n587), .A4(new_n588), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT113), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n950), .A2(new_n951), .A3(new_n956), .A4(KEYINPUT49), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n791), .A2(G1976), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n947), .A2(G8), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT52), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT112), .B(G1976), .Z(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n947), .A2(G8), .A3(new_n964), .A4(new_n960), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n959), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n945), .B2(new_n946), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT111), .B(new_n967), .C1(new_n945), .C2(new_n946), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n496), .B2(new_n508), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n942), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n970), .A2(new_n702), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT108), .B(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n942), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(G1971), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G303), .A2(G8), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(G8), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n966), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n487), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT71), .B1(new_n487), .B2(KEYINPUT4), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n494), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n504), .A2(new_n507), .ZN(new_n992));
  INV_X1    g567(.A(new_n501), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n944), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n972), .A2(new_n943), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n988), .B(new_n942), .C1(new_n998), .C2(new_n967), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n942), .A2(new_n967), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n947), .A2(KEYINPUT115), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n981), .B1(new_n1004), .B2(G2090), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n985), .B1(new_n1005), .B2(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n987), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1009));
  INV_X1    g584(.A(G2078), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n980), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n973), .B1(new_n968), .B2(new_n969), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n971), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(new_n751), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT45), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n942), .B1(new_n995), .B2(new_n1017), .ZN(new_n1018));
  OR4_X1    g593(.A1(new_n1015), .A2(new_n1016), .A3(G2078), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(G301), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1961), .B1(new_n1012), .B2(new_n971), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n509), .B2(new_n976), .ZN(new_n1022));
  NOR4_X1   g597(.A1(new_n978), .A2(new_n1022), .A3(new_n1015), .A4(G2078), .ZN(new_n1023));
  NOR4_X1   g598(.A1(new_n1021), .A2(new_n1011), .A3(new_n1023), .A4(G171), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1008), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1014), .A2(G301), .A3(new_n1019), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1021), .A2(new_n1011), .A3(new_n1023), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(KEYINPUT54), .C1(G301), .C2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1007), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n970), .A2(new_n1032), .A3(new_n971), .A4(new_n974), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1031), .B(G8), .C1(new_n1036), .C2(G286), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G168), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1040), .ZN(new_n1042));
  AOI211_X1 g617(.A(KEYINPUT123), .B(new_n1042), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1037), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g619(.A(new_n1031), .B(new_n1040), .C1(new_n1036), .C2(G8), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1030), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(new_n1038), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1036), .A2(G8), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT51), .A3(new_n1042), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(KEYINPUT124), .A3(new_n1050), .A4(new_n1037), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1029), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT56), .B(G2072), .Z(new_n1054));
  NOR3_X1   g629(.A1(new_n978), .A2(new_n979), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1956), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1004), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(G299), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n567), .A2(new_n575), .A3(KEYINPUT117), .A4(KEYINPUT57), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n569), .A2(new_n570), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n558), .B(new_n1062), .C1(new_n564), .C2(new_n566), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n1063), .B2(KEYINPUT57), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n567), .A2(new_n571), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1059), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1060), .A2(new_n1061), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1057), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n947), .A2(new_n1000), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1002), .B1(new_n1071), .B2(new_n988), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1956), .B1(new_n1072), .B2(new_n1001), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT118), .B(new_n1068), .C1(new_n1073), .C2(new_n1055), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1057), .B2(new_n1069), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n947), .A2(G2067), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1013), .B2(new_n734), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n877), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1053), .B(new_n1070), .C1(new_n1077), .C2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1055), .B(new_n1068), .C1(new_n1004), .C2(new_n1056), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1070), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1083), .B2(KEYINPUT122), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n877), .B1(new_n1079), .B2(KEYINPUT60), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1348), .B1(new_n1012), .B2(new_n971), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  NOR4_X1   g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n607), .A4(new_n1078), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1092), .A2(new_n1095), .B1(KEYINPUT60), .B2(new_n1079), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1057), .A2(new_n1069), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1083), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n980), .A2(new_n689), .ZN(new_n1100));
  INV_X1    g675(.A(new_n947), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT58), .B(G1341), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n548), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT59), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1096), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1091), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1052), .B1(new_n1085), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1046), .A2(new_n1051), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1007), .A2(new_n1020), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G288), .A2(G1976), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n959), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n951), .B(KEYINPUT114), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n949), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n966), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n986), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1007), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1036), .A2(G8), .A3(G168), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n985), .B1(new_n982), .B2(G8), .ZN(new_n1126));
  OR4_X1    g701(.A1(new_n1122), .A2(new_n987), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1121), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1109), .A2(new_n1115), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1022), .A2(new_n942), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n727), .B(G2067), .Z(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(G1996), .B2(new_n781), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n782), .A2(new_n689), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n811), .B(new_n815), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1137), .B(new_n1138), .C1(new_n819), .C2(new_n597), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n597), .A2(new_n819), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT109), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1131), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n781), .ZN(new_n1144));
  NOR2_X1   g719(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(G1996), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1131), .B1(new_n1133), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1130), .A2(G1996), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  AOI21_X1  g726(.A(new_n1130), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1141), .A2(KEYINPUT48), .A3(new_n1131), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT48), .B1(new_n1141), .B2(new_n1131), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n811), .A2(new_n814), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1136), .A2(new_n1156), .B1(G2067), .B2(new_n727), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1151), .B(new_n1155), .C1(new_n1131), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1143), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g734(.A(G319), .B1(new_n651), .B2(new_n652), .ZN(new_n1161));
  NOR2_X1   g735(.A1(G227), .A2(new_n1161), .ZN(new_n1162));
  AND3_X1   g736(.A1(new_n872), .A2(new_n696), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  AND3_X1   g738(.A1(new_n1163), .A2(new_n1164), .A3(new_n933), .ZN(new_n1165));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1163), .B2(new_n933), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1166), .ZN(G308));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n933), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n1168), .A2(KEYINPUT127), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n1163), .A2(new_n1164), .A3(new_n933), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1170), .ZN(G225));
endmodule


