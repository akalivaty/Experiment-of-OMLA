//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  OAI211_X1 g0045(.A(G1), .B(G13), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT65), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n248), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n255), .A2(G223), .B1(G77), .B2(new_n254), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n246), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n246), .A2(G274), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n245), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n246), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n215), .B2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G190), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(G200), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n209), .B1(new_n203), .B2(new_n244), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n273), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n210), .A2(G1), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(G50), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G50), .B2(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT9), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G58), .A2(G68), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n210), .B1(new_n288), .B2(new_n214), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n244), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n290), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n272), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n286), .A2(new_n287), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n287), .B1(new_n286), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n269), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n269), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n286), .A2(new_n297), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n266), .A2(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n266), .A2(G179), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n263), .B1(new_n312), .B2(new_n264), .ZN(new_n313));
  INV_X1    g0113(.A(G232), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n247), .B(new_n315), .C1(G226), .C2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n246), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n313), .A2(KEYINPUT13), .A3(new_n318), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n320), .A2(G179), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT70), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n320), .A2(new_n323), .A3(new_n321), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G169), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n326), .B2(KEYINPUT14), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(KEYINPUT14), .B2(new_n326), .ZN(new_n328));
  INV_X1    g0128(.A(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n279), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n329), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n214), .B2(new_n295), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n272), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT11), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n281), .A2(new_n329), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n334), .A2(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n331), .B(new_n338), .C1(new_n335), .C2(new_n334), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n324), .A2(G200), .A3(new_n325), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n267), .B1(new_n319), .B2(KEYINPUT13), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n339), .B1(new_n342), .B2(new_n321), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n222), .B2(new_n247), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G238), .B2(new_n255), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n263), .B1(new_n221), .B2(new_n264), .C1(new_n347), .C2(new_n246), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n350));
  OAI21_X1  g0150(.A(G190), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G200), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n290), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n292), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n270), .B1(new_n220), .B2(new_n279), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n336), .A2(G77), .A3(new_n282), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n351), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n349), .B2(new_n350), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n352), .A2(new_n307), .A3(new_n353), .ZN(new_n365));
  INV_X1    g0165(.A(new_n361), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n340), .A2(new_n344), .A3(new_n362), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n290), .A2(new_n281), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n280), .A2(new_n369), .B1(new_n279), .B2(new_n290), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(G58), .C2(G68), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n294), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n252), .A2(new_n253), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n251), .A2(KEYINPUT71), .A3(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT72), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT72), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT7), .A2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n383), .A2(new_n210), .A3(new_n384), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n329), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n392));
  AOI211_X1 g0192(.A(new_n373), .B(new_n381), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n247), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n329), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n373), .B1(new_n397), .B2(new_n381), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n270), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n372), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n270), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n254), .B2(new_n210), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n394), .B(G20), .C1(new_n252), .C2(new_n253), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n378), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n406), .B2(new_n373), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n387), .B1(new_n383), .B2(new_n384), .ZN(new_n409));
  INV_X1    g0209(.A(new_n389), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n391), .A2(KEYINPUT7), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  OAI211_X1 g0213(.A(KEYINPUT16), .B(new_n405), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n414), .A3(KEYINPUT74), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n371), .B1(new_n400), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n248), .B1(new_n383), .B2(new_n384), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n418));
  AND4_X1   g0218(.A1(KEYINPUT75), .A2(new_n385), .A3(G223), .A4(new_n248), .ZN(new_n419));
  AOI21_X1  g0219(.A(G1698), .B1(new_n383), .B2(new_n384), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT75), .B1(new_n420), .B2(G223), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n246), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n263), .B1(new_n314), .B2(new_n264), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n267), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(G200), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n416), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n416), .B2(new_n429), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT77), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n407), .A2(new_n414), .A3(KEYINPUT74), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT74), .B1(new_n407), .B2(new_n414), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n370), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n424), .A2(G179), .A3(new_n426), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n307), .B2(new_n428), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n438), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n433), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n428), .A2(G200), .ZN(new_n446));
  AOI211_X1 g0246(.A(G190), .B(new_n425), .C1(new_n422), .C2(new_n423), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n445), .B1(new_n438), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n416), .A2(new_n429), .A3(new_n431), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n435), .A2(new_n444), .A3(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n311), .A2(new_n368), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n273), .A2(G45), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n258), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n246), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(G257), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT79), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT4), .A2(G244), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n252), .A2(new_n253), .A3(new_n464), .A4(new_n248), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT78), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n247), .A2(new_n467), .A3(new_n248), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n252), .A2(new_n253), .A3(G250), .A4(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n221), .B1(new_n383), .B2(new_n384), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT4), .B1(new_n475), .B2(new_n248), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n463), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n385), .A2(G244), .A3(new_n248), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n472), .B1(new_n466), .B2(new_n468), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(KEYINPUT79), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT80), .B1(new_n483), .B2(new_n423), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n485), .B(new_n246), .C1(new_n477), .C2(new_n482), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n462), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G200), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  INV_X1    g0289(.A(G97), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n222), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n489), .B1(new_n493), .B2(KEYINPUT6), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n495));
  OAI21_X1  g0295(.A(G107), .B1(new_n402), .B2(new_n403), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n401), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n278), .A2(G97), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n273), .A2(G33), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n280), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n490), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n462), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n483), .B2(new_n423), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(G190), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n363), .B(new_n462), .C1(new_n484), .C2(new_n486), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n501), .A2(new_n490), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n507), .A2(new_n497), .A3(new_n498), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n474), .A2(new_n476), .A3(new_n463), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT79), .B1(new_n480), .B2(new_n481), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n423), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n462), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n512), .B2(new_n307), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n488), .A2(new_n505), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n420), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n385), .A2(G244), .A3(G1698), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n246), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n246), .A2(G274), .A3(new_n457), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n246), .A2(G250), .A3(new_n456), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT82), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n385), .A2(G238), .A3(new_n248), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n516), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n423), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n521), .A2(new_n522), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT82), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n307), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n524), .A2(new_n531), .A3(new_n363), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n385), .A2(new_n210), .A3(G68), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT19), .B1(new_n291), .B2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n210), .B1(new_n317), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n492), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n270), .B1(new_n279), .B2(new_n357), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n357), .B2(new_n501), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n533), .A2(new_n534), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n532), .A2(G200), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n524), .A2(new_n531), .A3(G190), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n543), .B1(new_n539), .B2(new_n501), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n280), .A2(G107), .A3(new_n500), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT86), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(KEYINPUT25), .C1(new_n278), .C2(G107), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT86), .B(KEYINPUT25), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n279), .A2(new_n222), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n210), .A2(G87), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT22), .B1(new_n247), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT84), .B1(new_n526), .B2(G20), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n210), .A3(G33), .A4(G116), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n222), .A3(G20), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n562), .A2(new_n564), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT22), .A2(G87), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n385), .A2(new_n210), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(new_n569), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n270), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT85), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n254), .B2(new_n559), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n580), .A3(new_n564), .ZN(new_n581));
  AOI211_X1 g0381(.A(G20), .B(new_n570), .C1(new_n383), .C2(new_n384), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT24), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n270), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n558), .B1(new_n577), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n420), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n385), .A2(G257), .A3(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n246), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n460), .A2(new_n223), .B1(new_n258), .B2(new_n458), .ZN(new_n592));
  OAI21_X1  g0392(.A(G169), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n385), .A2(G250), .A3(new_n248), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n423), .ZN(new_n598));
  INV_X1    g0398(.A(new_n592), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(G179), .A3(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n593), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n594), .B1(new_n593), .B2(new_n600), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n588), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n417), .A2(G264), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n385), .A2(G257), .A3(new_n248), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n254), .A2(G303), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n423), .ZN(new_n608));
  INV_X1    g0408(.A(new_n459), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n460), .A2(new_n217), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n608), .A2(G190), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n216), .B1(new_n273), .B2(G33), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n336), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n336), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n471), .B(new_n210), .C1(G33), .C2(new_n490), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n216), .A2(G20), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n270), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n619), .A2(new_n270), .A3(KEYINPUT20), .A4(new_n620), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n279), .B2(new_n216), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n459), .B(new_n610), .C1(new_n607), .C2(new_n423), .ZN(new_n628));
  INV_X1    g0428(.A(G200), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n612), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(G179), .A3(new_n626), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n307), .B1(new_n618), .B2(new_n625), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n630), .B(new_n631), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n558), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n586), .B1(new_n585), .B2(new_n270), .ZN(new_n639));
  AOI211_X1 g0439(.A(KEYINPUT85), .B(new_n401), .C1(new_n583), .C2(new_n584), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n629), .B1(new_n591), .B2(new_n592), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n598), .A2(new_n267), .A3(new_n599), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n603), .A2(new_n637), .A3(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n454), .A2(new_n514), .A3(new_n552), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n310), .ZN(new_n649));
  INV_X1    g0449(.A(new_n344), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n340), .B1(new_n650), .B2(new_n367), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n435), .A3(new_n452), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n444), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(new_n305), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n545), .A2(new_n550), .A3(new_n506), .A4(new_n513), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n506), .A2(new_n513), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n528), .A2(new_n529), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G200), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n547), .A2(new_n549), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n307), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n534), .A2(new_n544), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT26), .B1(new_n658), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n644), .B(new_n638), .C1(new_n640), .C2(new_n639), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n667), .A2(new_n663), .A3(new_n661), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n511), .A2(new_n485), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n483), .A2(KEYINPUT80), .A3(new_n423), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n503), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n505), .B1(new_n671), .B2(new_n629), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n610), .B1(new_n607), .B2(new_n423), .ZN(new_n673));
  AND4_X1   g0473(.A1(G179), .A2(new_n626), .A3(new_n673), .A4(new_n609), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n632), .A2(new_n633), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT21), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n593), .A2(new_n600), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n641), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n506), .A2(new_n513), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n668), .A2(new_n672), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n663), .B(KEYINPUT88), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n454), .B1(new_n666), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n654), .A2(new_n686), .ZN(G369));
  INV_X1    g0487(.A(new_n678), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n273), .A2(new_n210), .A3(G13), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n627), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT89), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n697), .B(KEYINPUT89), .C1(new_n637), .C2(new_n696), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n603), .A2(new_n646), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n588), .B2(new_n695), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n603), .A2(new_n694), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n678), .A2(new_n694), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n680), .B2(new_n694), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(G399));
  NOR2_X1   g0513(.A1(new_n540), .A2(G116), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  INV_X1    g0515(.A(new_n204), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n715), .A2(new_n273), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n208), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT28), .Z(new_n720));
  OAI21_X1  g0520(.A(new_n695), .B1(new_n666), .B2(new_n685), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT92), .B(new_n695), .C1(new_n666), .C2(new_n685), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n655), .A2(new_n656), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n658), .A2(new_n664), .A3(KEYINPUT26), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT94), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n656), .C1(new_n551), .C2(new_n682), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n602), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n641), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n678), .B1(new_n736), .B2(new_n601), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n668), .A3(new_n672), .A4(new_n682), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n684), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n694), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n723), .A2(KEYINPUT93), .A3(new_n724), .A4(new_n725), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n728), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT91), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n363), .B(new_n592), .C1(new_n597), .C2(new_n423), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n511), .A2(new_n462), .A3(new_n747), .A4(new_n673), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n748), .B2(new_n532), .ZN(new_n749));
  AOI21_X1  g0549(.A(G179), .B1(new_n598), .B2(new_n599), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n750), .A2(new_n632), .A3(new_n659), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n749), .A2(KEYINPUT30), .B1(new_n487), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n746), .B(new_n753), .C1(new_n748), .C2(new_n532), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n745), .B1(new_n755), .B2(new_n695), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n695), .B1(new_n752), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT31), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n647), .A2(new_n514), .A3(new_n552), .A4(new_n695), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G330), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n744), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n720), .B1(new_n763), .B2(G1), .ZN(G364));
  INV_X1    g0564(.A(G330), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n700), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT95), .Z(new_n767));
  AND2_X1   g0567(.A1(new_n210), .A2(G13), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n273), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n717), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n767), .A2(new_n702), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(G20), .B1(KEYINPUT96), .B2(G169), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(KEYINPUT96), .A2(G169), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n209), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n210), .A2(new_n363), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(G317), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n210), .A2(G190), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n363), .A3(new_n629), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OR3_X1    g0591(.A1(new_n629), .A2(KEYINPUT98), .A3(G179), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT98), .B1(new_n629), .B2(G179), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n210), .A2(new_n267), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n791), .A2(G329), .B1(G303), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n267), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n210), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n779), .A2(new_n267), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G294), .A2(new_n800), .B1(new_n801), .B2(G326), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n778), .A2(G190), .A3(new_n629), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n247), .B1(new_n804), .B2(G322), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G190), .A2(G200), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n778), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n792), .A2(new_n785), .A3(new_n793), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(G283), .B2(new_n811), .ZN(new_n812));
  AND4_X1   g0612(.A1(new_n784), .A2(new_n797), .A3(new_n802), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  OR3_X1    g0614(.A1(new_n786), .A2(KEYINPUT32), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n780), .ZN(new_n816));
  INV_X1    g0616(.A(new_n801), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n329), .C1(new_n214), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n808), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n254), .B1(new_n819), .B2(G77), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n800), .A2(G97), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n804), .A2(G58), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT32), .B1(new_n786), .B2(new_n814), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n795), .A2(new_n539), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n810), .A2(new_n222), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n818), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n777), .B1(new_n813), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n716), .A2(new_n254), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G355), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(G116), .B2(new_n204), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n386), .A2(new_n388), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n716), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n207), .A2(G45), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n242), .B2(G45), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(G13), .A2(G33), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(G20), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n777), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n771), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n828), .B1(new_n843), .B2(KEYINPUT97), .ZN(new_n844));
  INV_X1    g0644(.A(new_n839), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n701), .A2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(KEYINPUT97), .C2(new_n843), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n773), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n777), .A2(new_n837), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n772), .B1(new_n850), .B2(new_n220), .ZN(new_n851));
  INV_X1    g0651(.A(new_n777), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n790), .A2(new_n806), .B1(new_n539), .B2(new_n810), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  INV_X1    g0654(.A(G303), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n821), .B1(new_n816), .B2(new_n854), .C1(new_n855), .C2(new_n817), .ZN(new_n856));
  INV_X1    g0656(.A(G294), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n254), .B1(new_n808), .B2(new_n216), .C1(new_n857), .C2(new_n803), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n795), .A2(new_n222), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n853), .A2(new_n856), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n791), .A2(G132), .B1(G58), .B2(new_n800), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n810), .A2(new_n329), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G50), .B2(new_n796), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n861), .A2(new_n832), .A3(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n804), .A2(G143), .B1(new_n819), .B2(G159), .ZN(new_n865));
  INV_X1    g0665(.A(G137), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n865), .B1(new_n816), .B2(new_n293), .C1(new_n866), .C2(new_n817), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT34), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n860), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n367), .A2(new_n694), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n362), .B1(new_n361), .B2(new_n695), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n367), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n851), .B1(new_n852), .B2(new_n869), .C1(new_n872), .C2(new_n838), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n367), .ZN(new_n874));
  INV_X1    g0674(.A(new_n870), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n723), .A2(new_n725), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n872), .B(new_n695), .C1(new_n666), .C2(new_n685), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n762), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT100), .A3(new_n772), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n762), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT100), .B1(new_n879), .B2(new_n772), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(G384));
  OR2_X1    g0684(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n211), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  AND4_X1   g0688(.A1(G77), .A2(new_n208), .A3(new_n376), .A4(new_n377), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n889), .A2(KEYINPUT101), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n889), .A2(KEYINPUT101), .B1(new_n214), .B2(G68), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n273), .B(G13), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n728), .A2(new_n454), .A3(new_n742), .A4(new_n743), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n654), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n381), .B1(new_n390), .B2(new_n392), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n373), .A2(KEYINPUT103), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n272), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n692), .B1(new_n900), .B2(new_n370), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n453), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n370), .ZN(new_n903));
  INV_X1    g0703(.A(new_n692), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n441), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n416), .A2(new_n429), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n438), .A2(new_n441), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n438), .A2(new_n904), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(new_n906), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(KEYINPUT37), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n911), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n449), .A2(new_n451), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n444), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n914), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n340), .A2(new_n694), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n902), .A2(new_n912), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n914), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n913), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n922), .B(new_n923), .C1(new_n926), .C2(new_n921), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n339), .A2(new_n694), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n340), .A2(new_n344), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n339), .B(new_n694), .C1(new_n328), .C2(new_n650), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n878), .A2(KEYINPUT102), .A3(new_n875), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT102), .B1(new_n878), .B2(new_n875), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n926), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n692), .B1(new_n442), .B2(new_n443), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n927), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n895), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n759), .B1(KEYINPUT31), .B2(new_n757), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n757), .A2(KEYINPUT31), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT104), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n876), .B1(new_n929), .B2(new_n930), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT104), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n756), .A2(new_n943), .A3(new_n758), .A4(new_n759), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT40), .B1(new_n925), .B2(new_n913), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n913), .A2(new_n919), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT40), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n941), .A2(new_n944), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n454), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n765), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n951), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n938), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n273), .B2(new_n768), .C1(new_n938), .C2(new_n955), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n893), .B1(new_n958), .B2(new_n959), .ZN(G367));
  NAND2_X1  g0760(.A1(new_n502), .A2(new_n694), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n514), .A2(new_n961), .B1(new_n658), .B2(new_n694), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n710), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n672), .A2(new_n603), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n694), .B1(new_n966), .B2(new_n682), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n964), .B2(KEYINPUT42), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n548), .A2(new_n694), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n684), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n664), .B2(new_n969), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n965), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n708), .A2(new_n962), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n975), .B(new_n976), .Z(new_n977));
  XOR2_X1   g0777(.A(new_n717), .B(KEYINPUT41), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n711), .A2(new_n962), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT44), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n711), .A2(new_n962), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n708), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n707), .A2(new_n709), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(new_n702), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n763), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n978), .B1(new_n990), .B2(new_n763), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n977), .B1(new_n991), .B2(new_n770), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n840), .B1(new_n204), .B2(new_n357), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n833), .B2(new_n235), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n772), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G107), .A2(new_n800), .B1(new_n801), .B2(G311), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n857), .B2(new_n816), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n810), .A2(new_n490), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G303), .A2(new_n804), .B1(new_n787), .B2(G317), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n854), .B2(new_n808), .ZN(new_n1000));
  OR4_X1    g0800(.A1(new_n832), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n795), .A2(new_n216), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT46), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n799), .A2(new_n329), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G143), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n816), .B2(new_n814), .C1(new_n1006), .C2(new_n817), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n803), .A2(new_n293), .B1(new_n808), .B2(new_n214), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n254), .B(new_n1008), .C1(G137), .C2(new_n787), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n796), .A2(G58), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n220), .C2(new_n810), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1001), .A2(new_n1003), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n995), .B1(new_n852), .B2(new_n1013), .C1(new_n972), .C2(new_n845), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n992), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n763), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n989), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n717), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1018), .A2(KEYINPUT108), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(KEYINPUT108), .B2(new_n1018), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n705), .A2(new_n706), .A3(new_n839), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n799), .A2(new_n357), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n814), .B2(new_n817), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n355), .B2(new_n780), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n803), .A2(new_n214), .B1(new_n808), .B2(new_n329), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1026), .B(new_n998), .C1(G150), .C2(new_n787), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n796), .A2(G77), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n832), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n832), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n811), .A2(G116), .B1(G326), .B2(new_n787), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n795), .A2(new_n857), .B1(new_n854), .B2(new_n799), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n804), .A2(G317), .B1(new_n819), .B2(G303), .ZN(new_n1033));
  INV_X1    g0833(.A(G322), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(new_n816), .B2(new_n806), .C1(new_n1034), .C2(new_n817), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1030), .B(new_n1031), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1029), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n777), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n232), .A2(new_n259), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1044), .A2(new_n833), .B1(new_n715), .B2(new_n829), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n290), .A2(G50), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT50), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n259), .B1(new_n329), .B2(new_n220), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n715), .B(new_n1048), .C1(new_n1047), .C2(new_n1046), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1045), .A2(new_n1049), .B1(G107), .B2(new_n204), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n772), .B1(new_n1050), .B2(new_n840), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1051), .B2(KEYINPUT107), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(KEYINPUT107), .B2(new_n1051), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n989), .A2(new_n770), .B1(new_n1021), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1020), .A2(new_n1054), .ZN(G393));
  OAI22_X1  g0855(.A1(new_n817), .A2(new_n293), .B1(new_n814), .B2(new_n803), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT51), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n799), .A2(new_n220), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1006), .A2(new_n786), .B1(new_n808), .B2(new_n290), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G50), .C2(new_n780), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G68), .A2(new_n796), .B1(new_n811), .B2(G87), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n832), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT109), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n816), .A2(new_n855), .B1(new_n216), .B2(new_n799), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT110), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n817), .A2(new_n781), .B1(new_n806), .B2(new_n803), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n254), .B1(new_n808), .B2(new_n857), .C1(new_n1034), .C2(new_n786), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n826), .B(new_n1068), .C1(G283), .C2(new_n796), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1063), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1062), .A2(KEYINPUT109), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n777), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n833), .A2(new_n239), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n841), .B1(G97), .B2(new_n716), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n772), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n962), .B2(new_n839), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n984), .B2(new_n770), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n990), .A2(new_n717), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n984), .B1(new_n763), .B2(new_n989), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(G390));
  NAND4_X1  g0882(.A1(new_n941), .A2(new_n942), .A3(new_n944), .A4(G330), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT112), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n922), .B1(new_n926), .B2(new_n921), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n878), .A2(new_n875), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT102), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n878), .A2(KEYINPUT102), .A3(new_n875), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n931), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1087), .B1(new_n1092), .B2(new_n923), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n733), .A2(new_n731), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n732), .B1(new_n655), .B2(new_n656), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n695), .B(new_n874), .C1(new_n1096), .C2(new_n739), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n931), .B1(new_n1097), .B2(new_n875), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n923), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n920), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT111), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT111), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n923), .B1(new_n913), .B2(new_n919), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n870), .B1(new_n741), .B2(new_n874), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1103), .C1(new_n1104), .C2(new_n931), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1086), .B1(new_n1093), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(G330), .B(new_n872), .C1(new_n939), .C2(new_n940), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1109), .A2(new_n931), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1093), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n952), .A2(G330), .A3(new_n454), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n894), .A2(new_n654), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n941), .A2(G330), .A3(new_n944), .A4(new_n872), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n931), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1110), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1104), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1109), .A2(new_n931), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1083), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT113), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT113), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1119), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1108), .A2(new_n1112), .A3(new_n1115), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1115), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1099), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1130), .A2(new_n1087), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1112), .B1(new_n1131), .B2(new_n1086), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1127), .A2(new_n1133), .A3(new_n717), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1112), .B(new_n770), .C1(new_n1131), .C2(new_n1086), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n850), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n817), .A2(new_n854), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1058), .B(new_n1137), .C1(G107), .C2(new_n780), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n247), .B1(new_n804), .B2(G116), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n539), .B2(new_n795), .C1(new_n490), .C2(new_n808), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n862), .B(new_n1140), .C1(G294), .C2(new_n791), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n247), .B1(new_n808), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G132), .B2(new_n804), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n214), .B2(new_n810), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G159), .A2(new_n800), .B1(new_n780), .B2(G137), .ZN(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n817), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1145), .B(new_n1148), .C1(G125), .C2(new_n791), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n795), .A2(new_n293), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1138), .A2(new_n1141), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n771), .B1(new_n355), .B2(new_n1136), .C1(new_n1153), .C2(new_n852), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1087), .B2(new_n837), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT115), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT116), .B1(new_n1135), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1135), .A2(KEYINPUT116), .A3(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1134), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1134), .B(KEYINPUT117), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(G378));
  INV_X1    g0963(.A(KEYINPUT55), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n306), .B2(new_n904), .ZN(new_n1165));
  AOI211_X1 g0965(.A(KEYINPUT55), .B(new_n692), .C1(new_n286), .C2(new_n297), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n311), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n305), .A2(new_n310), .A3(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1169), .B1(new_n305), .B2(new_n310), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n649), .B(new_n1167), .C1(new_n302), .C2(new_n304), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n837), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1005), .B1(new_n222), .B2(new_n803), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n811), .A2(G58), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1028), .B(new_n1180), .C1(new_n790), .C2(new_n854), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G116), .C2(new_n801), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n816), .A2(new_n490), .B1(new_n357), .B2(new_n808), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT118), .Z(new_n1184));
  NAND4_X1  g0984(.A1(new_n1182), .A2(new_n245), .A3(new_n1030), .A4(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT58), .Z(new_n1186));
  OAI22_X1  g0986(.A1(new_n803), .A2(new_n1147), .B1(new_n808), .B2(new_n866), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G132), .B2(new_n780), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G150), .A2(new_n800), .B1(new_n801), .B2(G125), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n795), .C2(new_n1142), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n811), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G50), .B1(new_n244), .B2(new_n245), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n832), .B2(G41), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n777), .B1(new_n1186), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n772), .B1(new_n850), .B2(new_n214), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1178), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n920), .A2(new_n941), .A3(new_n944), .A4(new_n942), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(KEYINPUT40), .A2(new_n1204), .B1(new_n945), .B2(new_n946), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1177), .B1(new_n1205), .B2(new_n765), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n937), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1177), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n951), .A2(G330), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT122), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1206), .A2(new_n1209), .A3(new_n1207), .A4(KEYINPUT122), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1208), .B1(new_n951), .B2(G330), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n765), .B(new_n1177), .C1(new_n947), .C2(new_n950), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n937), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT121), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1207), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT121), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1214), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1203), .B1(new_n1222), .B2(new_n770), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT123), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1093), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n1107), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1114), .B1(new_n1226), .B2(new_n1126), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1219), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1224), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1217), .B2(new_n1210), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1119), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1125), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n1123), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1115), .B1(new_n1132), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1232), .A2(new_n1236), .A3(KEYINPUT123), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1230), .A2(new_n717), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1236), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1223), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT124), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(KEYINPUT124), .B(new_n1223), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(G375));
  NAND2_X1  g1045(.A1(new_n931), .A2(new_n837), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n771), .B1(new_n1136), .B2(G68), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n791), .A2(G128), .B1(G159), .B2(new_n796), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n800), .A2(G50), .B1(new_n819), .B2(G150), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n832), .A3(new_n1180), .A4(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT127), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n801), .A2(G132), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1252), .B1(new_n866), .B2(new_n803), .C1(new_n816), .C2(new_n1142), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT126), .Z(new_n1254));
  OAI22_X1  g1054(.A1(new_n790), .A2(new_n855), .B1(new_n490), .B2(new_n795), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT125), .Z(new_n1256));
  OAI221_X1 g1056(.A(new_n1023), .B1(new_n816), .B2(new_n216), .C1(new_n857), .C2(new_n817), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n810), .A2(new_n220), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n254), .B1(new_n808), .B2(new_n222), .C1(new_n854), .C2(new_n803), .ZN(new_n1259));
  OR3_X1    g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1251), .A2(new_n1254), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1247), .B1(new_n1261), .B2(new_n777), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1126), .A2(new_n770), .B1(new_n1246), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n978), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1128), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1126), .A2(new_n1115), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1263), .B1(new_n1265), .B2(new_n1266), .ZN(G381));
  NOR4_X1   g1067(.A1(G387), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1159), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1244), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n693), .A2(G213), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1244), .A2(new_n1269), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(G213), .A3(new_n1274), .ZN(G409));
  NAND3_X1  g1075(.A1(new_n1222), .A2(new_n1264), .A3(new_n1236), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1217), .A2(new_n1210), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1203), .B1(new_n1277), .B2(new_n770), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1269), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1240), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1266), .B1(KEYINPUT60), .B2(new_n1128), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1235), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n717), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1263), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(G384), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G384), .B(new_n1263), .C1(new_n1283), .C2(new_n1285), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1282), .A2(new_n1272), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1273), .A2(G2897), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1290), .B(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1159), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1222), .A2(new_n770), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1202), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1232), .A2(new_n1236), .A3(KEYINPUT123), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT123), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n717), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1222), .A2(new_n1236), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1231), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1299), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1297), .B1(new_n1306), .B2(G378), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1296), .B1(new_n1307), .B2(new_n1273), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1282), .A2(new_n1309), .A3(new_n1272), .A4(new_n1291), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1293), .A2(new_n1294), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(G390), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G387), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n848), .B1(new_n1020), .B2(new_n1054), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(G387), .A2(new_n1312), .ZN(new_n1316));
  OR4_X1    g1116(.A1(new_n1270), .A2(new_n1314), .A3(new_n1315), .A4(new_n1316), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1270), .A2(new_n1315), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1319), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1282), .A2(new_n1272), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1296), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1292), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1282), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1291), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1321), .A2(new_n1323), .A3(new_n1325), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1327), .ZN(G405));
  NAND3_X1  g1128(.A1(new_n1242), .A2(new_n1269), .A3(new_n1243), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1306), .A2(G378), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1290), .A3(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1290), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1319), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1333), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1321), .A3(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(G402));
endmodule


