//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n533, new_n534, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT68), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT69), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT70), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT71), .ZN(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(G136), .B2(new_n465), .ZN(G162));
  AND2_X1   g054(.A1(KEYINPUT72), .A2(G138), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n466), .B(new_n480), .C1(new_n462), .C2(new_n463), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT4), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n474), .B2(G126), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G164));
  NAND2_X1  g063(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n489));
  INV_X1    g064(.A(G543), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n493), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT6), .B(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G50), .ZN(new_n499));
  AND3_X1   g074(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(G543), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT74), .B(G88), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n498), .A2(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n496), .A2(new_n506), .ZN(G166));
  XOR2_X1   g082(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n508));
  NAND3_X1  g083(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n493), .A2(G63), .A3(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n498), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G51), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n504), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G89), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(G168));
  AOI22_X1  g092(.A1(new_n493), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n495), .ZN(new_n519));
  INV_X1    g094(.A(G52), .ZN(new_n520));
  INV_X1    g095(.A(G90), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n498), .A2(new_n520), .B1(new_n504), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G171));
  OAI211_X1 g098(.A(G43), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n524));
  INV_X1    g099(.A(G81), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n504), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(G56), .B1(new_n500), .B2(new_n501), .ZN(new_n527));
  NAND2_X1  g102(.A1(G68), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n495), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G860), .ZN(G153));
  NAND4_X1  g106(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g107(.A1(G1), .A2(G3), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT8), .ZN(new_n534));
  NAND4_X1  g109(.A1(G319), .A2(G483), .A3(G661), .A4(new_n534), .ZN(G188));
  OAI211_X1 g110(.A(G53), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT9), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT9), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n497), .A2(new_n538), .A3(G53), .A4(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(G91), .ZN(new_n541));
  INV_X1    g116(.A(G65), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n491), .B2(new_n492), .ZN(new_n543));
  AND2_X1   g118(.A1(G78), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n540), .A2(new_n541), .A3(new_n548), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G299));
  INV_X1    g126(.A(G171), .ZN(G301));
  INV_X1    g127(.A(G168), .ZN(G286));
  INV_X1    g128(.A(G166), .ZN(G303));
  NAND2_X1  g129(.A1(new_n512), .A2(G49), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n515), .A2(G87), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n493), .B2(G74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(G288));
  AOI22_X1  g133(.A1(new_n493), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n495), .ZN(new_n560));
  INV_X1    g135(.A(G48), .ZN(new_n561));
  INV_X1    g136(.A(G86), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n498), .A2(new_n561), .B1(new_n504), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G305));
  AOI22_X1  g140(.A1(new_n493), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n495), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G47), .ZN(new_n569));
  INV_X1    g144(.A(G85), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n498), .A2(new_n569), .B1(new_n504), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n568), .A2(new_n571), .ZN(G290));
  NAND2_X1  g147(.A1(G301), .A2(G868), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n493), .A2(G66), .ZN(new_n574));
  NAND2_X1  g149(.A1(G79), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n579), .A3(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  INV_X1    g157(.A(G92), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n504), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n581), .A2(new_n584), .B1(G54), .B2(new_n512), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n573), .B1(new_n587), .B2(G868), .ZN(G321));
  XOR2_X1   g163(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G868), .B2(new_n550), .ZN(G297));
  OAI21_X1  g166(.A(new_n590), .B1(G868), .B2(new_n550), .ZN(G280));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n587), .B1(new_n593), .B2(G860), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT79), .Z(G148));
  NAND3_X1  g170(.A1(new_n493), .A2(G81), .A3(new_n497), .ZN(new_n596));
  INV_X1    g171(.A(new_n528), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n493), .B2(G56), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n524), .B(new_n596), .C1(new_n598), .C2(new_n495), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n587), .A2(KEYINPUT80), .A3(new_n593), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n586), .B2(G559), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  MUX2_X1   g178(.A(new_n599), .B(new_n603), .S(G868), .Z(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g180(.A(new_n464), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n467), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n465), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n474), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n466), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT84), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n632), .B(new_n633), .Z(new_n634));
  OR2_X1    g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT18), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n648), .A2(new_n643), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n644), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n643), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n647), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT87), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n662), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G27), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G164), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT98), .ZN(new_n682));
  INV_X1    g257(.A(G2078), .ZN(new_n683));
  NOR2_X1   g258(.A1(G4), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n587), .B2(G16), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n682), .A2(new_n683), .B1(G1348), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(G1348), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n687), .C1(new_n683), .C2(new_n682), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT90), .B(G16), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G20), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n550), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1956), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G171), .A2(new_n693), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G5), .B2(new_n693), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n679), .A2(G33), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n465), .A2(G139), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n606), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(new_n466), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n472), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G34), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n679), .B1(new_n712), .B2(G34), .ZN(new_n714));
  OAI22_X1  g289(.A1(new_n711), .A2(new_n679), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G162), .A2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G29), .B2(G35), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT29), .B(G2090), .Z(new_n720));
  AOI211_X1 g295(.A(new_n710), .B(new_n717), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n693), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n693), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n719), .A2(new_n720), .ZN(new_n726));
  INV_X1    g301(.A(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n729));
  OR2_X1    g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n617), .B2(new_n679), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n708), .A2(new_n709), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n726), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND4_X1   g310(.A1(new_n700), .A2(new_n721), .A3(new_n725), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n679), .A2(G26), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(G128), .A2(new_n474), .B1(new_n465), .B2(G140), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  INV_X1    g316(.A(G116), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(G2067), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(G2067), .ZN(new_n749));
  INV_X1    g324(.A(new_n689), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G19), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n530), .B2(new_n750), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1341), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n748), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n698), .A2(new_n699), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT97), .Z(new_n756));
  AND2_X1   g331(.A1(new_n679), .A2(G32), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n474), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n696), .A2(new_n736), .A3(new_n754), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G6), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n564), .B2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT32), .B(G1981), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n750), .A2(G22), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n750), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n693), .A2(G23), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n555), .A2(new_n557), .A3(new_n556), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n693), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n776), .A2(new_n777), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n679), .A2(G25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n465), .A2(G131), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n474), .A2(G119), .ZN(new_n792));
  OR2_X1    g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(new_n679), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  XOR2_X1   g374(.A(new_n798), .B(new_n799), .Z(new_n800));
  NOR2_X1   g375(.A1(new_n750), .A2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G290), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n750), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1986), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n788), .A2(new_n789), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT36), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n788), .A2(new_n808), .A3(new_n789), .A4(new_n805), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n770), .B1(new_n807), .B2(new_n809), .ZN(G311));
  XNOR2_X1  g385(.A(G311), .B(KEYINPUT100), .ZN(G150));
  OAI211_X1 g386(.A(G55), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n504), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(G67), .B1(new_n500), .B2(new_n501), .ZN(new_n815));
  NAND2_X1  g390(.A1(G80), .A2(G543), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n495), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT105), .B(G860), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n493), .A2(G93), .A3(new_n497), .ZN(new_n822));
  INV_X1    g397(.A(new_n816), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n493), .B2(G67), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n812), .B(new_n822), .C1(new_n824), .C2(new_n495), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT102), .B1(new_n530), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n530), .A2(new_n825), .A3(KEYINPUT102), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n818), .A2(new_n599), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(new_n818), .B2(new_n599), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n826), .A2(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT104), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n587), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n819), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n821), .B1(new_n838), .B2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n617), .B(new_n711), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(G162), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n765), .B(G164), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(new_n795), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n795), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(G130), .A2(new_n474), .B1(new_n465), .B2(G142), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n848), .A2(new_n466), .A3(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n466), .B2(G118), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT107), .ZN(new_n853));
  INV_X1    g428(.A(new_n608), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(new_n745), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n707), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n846), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n846), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n842), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  INV_X1    g441(.A(new_n842), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n862), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g446(.A(KEYINPUT110), .ZN(new_n872));
  XNOR2_X1  g447(.A(G288), .B(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(new_n564), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n564), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(G303), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(G290), .B(G166), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n874), .B2(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT42), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n600), .A2(new_n884), .A3(new_n602), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n600), .B2(new_n602), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n831), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n603), .A2(KEYINPUT108), .ZN(new_n889));
  INV_X1    g464(.A(new_n831), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n547), .A2(new_n585), .A3(new_n549), .A4(new_n580), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n547), .A2(new_n549), .B1(new_n580), .B2(new_n585), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n550), .A2(new_n586), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(KEYINPUT41), .A3(new_n894), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n899), .A3(KEYINPUT109), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n893), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n881), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n888), .A2(new_n891), .A3(new_n901), .ZN(new_n908));
  AND4_X1   g483(.A1(new_n883), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n883), .A2(new_n907), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n818), .A2(G868), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n883), .A2(new_n907), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n905), .A2(new_n908), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n883), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI211_X1 g494(.A(KEYINPUT111), .B(new_n912), .C1(new_n919), .C2(G868), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n911), .B2(new_n913), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n818), .B2(new_n599), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n530), .A2(new_n825), .A3(KEYINPUT102), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n530), .B2(new_n825), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n818), .A2(new_n599), .A3(new_n828), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n928), .A2(new_n931), .A3(G301), .ZN(new_n932));
  AOI21_X1  g507(.A(G301), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(G286), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n831), .A2(G171), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n928), .A2(new_n931), .A3(G301), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(G168), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n937), .A3(new_n901), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n934), .A2(new_n937), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n897), .A2(new_n899), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n941), .B2(new_n882), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n932), .A2(new_n933), .A3(G286), .ZN(new_n944));
  AOI21_X1  g519(.A(G168), .B1(new_n935), .B2(new_n936), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n903), .B(new_n900), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n881), .A3(new_n938), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n900), .A2(new_n903), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n938), .B1(new_n939), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n882), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(KEYINPUT112), .A3(new_n869), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n881), .B1(new_n946), .B2(new_n938), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(G37), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n949), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n924), .B(new_n948), .C1(new_n957), .C2(new_n943), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n947), .A2(new_n943), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n953), .B2(new_n956), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n943), .B1(new_n942), .B2(new_n947), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  AOI21_X1  g538(.A(G1384), .B1(new_n482), .B2(new_n486), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n965), .A2(KEYINPUT113), .ZN(new_n966));
  XOR2_X1   g541(.A(KEYINPUT114), .B(G40), .Z(new_n967));
  AND3_X1   g542(.A1(new_n468), .A2(new_n472), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n965), .B2(KEYINPUT113), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1986), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n802), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(G1986), .A3(G290), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT115), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n765), .A2(G1996), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n765), .A2(G1996), .ZN(new_n978));
  INV_X1    g553(.A(G2067), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n745), .B(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n971), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n971), .A3(KEYINPUT116), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n795), .B(new_n799), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n984), .B(new_n985), .C1(new_n970), .C2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n976), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n968), .A2(new_n964), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n783), .A2(G1976), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(G8), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n783), .A2(G1976), .ZN(new_n992));
  OR3_X1    g567(.A1(new_n991), .A2(KEYINPUT52), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(KEYINPUT52), .ZN(new_n994));
  OR3_X1    g569(.A1(new_n560), .A2(new_n563), .A3(G1981), .ZN(new_n995));
  OAI21_X1  g570(.A(G1981), .B1(new_n560), .B2(new_n563), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(KEYINPUT119), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n998));
  NAND3_X1  g573(.A1(G305), .A2(new_n998), .A3(G1981), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n989), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n997), .B2(new_n999), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n993), .B(new_n994), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n968), .B1(new_n964), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT118), .B1(new_n964), .B2(new_n1008), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n964), .A2(KEYINPUT118), .A3(new_n1008), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2090), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n968), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(new_n1017), .A3(KEYINPUT117), .A4(new_n968), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1022), .A3(new_n780), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1003), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G166), .A2(new_n1003), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT55), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1007), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1009), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n964), .A2(new_n1008), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1014), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1023), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1026), .B1(new_n1031), .B2(G8), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1021), .A2(new_n1017), .A3(new_n968), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1013), .A2(new_n716), .B1(new_n724), .B2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(new_n1003), .A3(G286), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1027), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT63), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1026), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1027), .A2(new_n1043), .A3(KEYINPUT63), .A4(new_n1036), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1046));
  INV_X1    g621(.A(G1956), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n546), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT121), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n541), .A2(new_n545), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT120), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n540), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1052), .A2(KEYINPUT120), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1049), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1048), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1057), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1002), .A2(new_n979), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1013), .B2(G1348), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n587), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1012), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1028), .B1(new_n1069), .B2(new_n1010), .ZN(new_n1070));
  INV_X1    g645(.A(G1348), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1070), .A2(new_n1071), .B1(new_n979), .B2(new_n1002), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n586), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n989), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n989), .A2(KEYINPUT122), .A3(new_n1074), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1077), .B(new_n1078), .C1(new_n1034), .C2(G1996), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n530), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1079), .B2(new_n530), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n586), .A2(KEYINPUT123), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT60), .B1(new_n586), .B2(KEYINPUT123), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1066), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1072), .A2(KEYINPUT60), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1064), .A2(new_n1090), .A3(new_n1061), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT61), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1068), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1070), .A2(G2084), .B1(G1966), .B2(new_n1058), .ZN(new_n1096));
  OAI21_X1  g671(.A(G8), .B1(new_n1096), .B2(G286), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1035), .A2(G168), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT51), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1003), .B1(new_n1035), .B2(G168), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n966), .A2(new_n969), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G160), .A2(G40), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT124), .ZN(new_n1106));
  NAND2_X1  g681(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1107));
  OR2_X1    g682(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1108));
  AND4_X1   g683(.A1(KEYINPUT53), .A2(new_n1017), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1070), .A2(new_n699), .ZN(new_n1111));
  AOI21_X1  g686(.A(G2078), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1110), .B(new_n1111), .C1(new_n1112), .C2(KEYINPUT53), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G171), .B(KEYINPUT54), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1058), .A2(KEYINPUT53), .A3(new_n683), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1111), .B(new_n1116), .C1(new_n1112), .C2(KEYINPUT53), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1114), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1095), .A2(new_n1103), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1045), .B1(new_n1094), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1096), .A2(G286), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1101), .B1(new_n1100), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT62), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1099), .A2(new_n1125), .A3(new_n1102), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1117), .A2(G171), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1124), .A2(new_n1126), .A3(new_n1095), .A4(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1041), .A2(new_n1007), .A3(new_n1042), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n995), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1132), .B2(new_n1004), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n988), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n973), .B(KEYINPUT48), .Z(new_n1136));
  INV_X1    g711(.A(new_n765), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n970), .B1(new_n1137), .B2(new_n980), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n970), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT46), .B1(new_n970), .B2(G1996), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT47), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n987), .A2(new_n1136), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n984), .A2(new_n797), .A3(new_n799), .A4(new_n985), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(G2067), .B2(new_n745), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n970), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1135), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g727(.A(new_n948), .B1(new_n957), .B2(new_n943), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n658), .A2(G319), .ZN(new_n1155));
  AOI21_X1  g729(.A(new_n1155), .B1(new_n639), .B2(new_n640), .ZN(new_n1156));
  OAI21_X1  g730(.A(new_n677), .B1(KEYINPUT127), .B2(new_n1156), .ZN(new_n1157));
  AND2_X1   g731(.A1(new_n1156), .A2(KEYINPUT127), .ZN(new_n1158));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g733(.A1(new_n1154), .A2(new_n1159), .A3(new_n870), .ZN(G308));
  NAND3_X1  g734(.A1(new_n1154), .A2(new_n1159), .A3(new_n870), .ZN(G225));
endmodule


