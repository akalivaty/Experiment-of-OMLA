//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(G128), .B(new_n189), .C1(new_n190), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n195), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n193), .A2(new_n206), .A3(new_n209), .A4(new_n197), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n215), .A2(KEYINPUT11), .B1(new_n216), .B2(G137), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT64), .A4(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n215), .A2(KEYINPUT11), .B1(new_n216), .B2(G137), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n214), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AND4_X1   g038(.A1(KEYINPUT64), .A2(new_n218), .A3(new_n219), .A4(G134), .ZN(new_n225));
  AOI22_X1  g039(.A1(KEYINPUT64), .A2(new_n218), .B1(new_n219), .B2(G134), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n214), .B(new_n222), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n213), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n228), .A3(KEYINPUT12), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G101), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n234), .A2(KEYINPUT75), .A3(new_n235), .A4(G101), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT0), .A4(G128), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n194), .A2(new_n195), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT0), .B(G128), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n234), .B2(G101), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n206), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT10), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n240), .A2(new_n246), .B1(new_n247), .B2(new_n212), .ZN(new_n248));
  INV_X1    g062(.A(new_n228), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n210), .A2(KEYINPUT76), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n193), .A2(new_n197), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n206), .A2(new_n209), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT10), .A4(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n249), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n233), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(G110), .B(G140), .Z(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT74), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n259), .A2(G227), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n240), .A2(new_n246), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n212), .A2(new_n247), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n254), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n228), .ZN(new_n266));
  INV_X1    g080(.A(new_n261), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n255), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G469), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  INV_X1    g086(.A(new_n268), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n267), .B1(new_n233), .B2(new_n255), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT77), .A3(G469), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n233), .A2(new_n255), .A3(new_n267), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n267), .B1(new_n266), .B2(new_n255), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n270), .B(new_n272), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G214), .B1(G237), .B2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G125), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n193), .A2(new_n283), .A3(new_n197), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n241), .B(G125), .C1(new_n242), .C2(new_n243), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n259), .A2(G224), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n284), .A2(new_n285), .A3(new_n288), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n250), .A2(new_n253), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G116), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G119), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT2), .B(G113), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G116), .B(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT5), .ZN(new_n303));
  OAI21_X1  g117(.A(G113), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n299), .A2(new_n300), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT2), .B(G113), .Z(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n302), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n245), .A2(new_n206), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n294), .A2(new_n306), .B1(new_n240), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G122), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n293), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n304), .B1(new_n303), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n302), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n301), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n210), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n312), .B(KEYINPUT8), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n305), .A2(new_n303), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n309), .ZN(new_n322));
  INV_X1    g136(.A(new_n210), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n314), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n312), .B(KEYINPUT8), .Z(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n306), .B2(new_n210), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(KEYINPUT80), .C1(new_n210), .C2(new_n318), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G902), .B1(new_n313), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n240), .A2(new_n310), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n306), .A2(new_n250), .A3(new_n253), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n312), .A2(KEYINPUT6), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n335), .ZN(new_n337));
  AOI211_X1 g151(.A(KEYINPUT78), .B(new_n337), .C1(new_n332), .C2(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(new_n333), .A3(new_n312), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT6), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n312), .B1(new_n332), .B2(new_n333), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n336), .A2(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n284), .A2(new_n285), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n286), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n330), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT82), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n312), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n334), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n339), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n352), .B(new_n344), .C1(new_n338), .C2(new_n336), .ZN(new_n353));
  INV_X1    g167(.A(new_n348), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n330), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n282), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT72), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n272), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G221), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n360), .B(KEYINPUT73), .Z(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n283), .A2(G140), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT70), .A4(KEYINPUT16), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT16), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT16), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n363), .A3(G125), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT70), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n191), .B(new_n366), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n364), .A2(new_n365), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n370), .B(new_n369), .C1(new_n374), .C2(new_n368), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n191), .B1(new_n375), .B2(new_n366), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(G237), .A2(G953), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(G143), .A3(G214), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n378), .B2(G214), .ZN(new_n381));
  OAI21_X1  g195(.A(G131), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT84), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n259), .A3(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n188), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n379), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n214), .A3(new_n379), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n383), .A2(new_n384), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n388), .B2(G131), .ZN(new_n393));
  AOI211_X1 g207(.A(KEYINPUT84), .B(new_n214), .C1(new_n387), .C2(new_n379), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT17), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n377), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n374), .A2(G146), .ZN(new_n398));
  XNOR2_X1  g212(.A(G125), .B(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n191), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n387), .A2(new_n379), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(G113), .B(G122), .Z(new_n406));
  XOR2_X1   g220(.A(KEYINPUT86), .B(G104), .Z(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT87), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n404), .A4(new_n408), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n272), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G475), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n404), .A2(new_n408), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n399), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n374), .B1(new_n419), .B2(KEYINPUT19), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(G146), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n376), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n415), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n408), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n405), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n414), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n408), .B1(new_n396), .B2(new_n404), .ZN(new_n429));
  INV_X1    g243(.A(new_n427), .ZN(new_n430));
  NOR4_X1   g244(.A1(new_n429), .A2(new_n424), .A3(KEYINPUT20), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n413), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G128), .B(G143), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n216), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n297), .B2(G122), .ZN(new_n436));
  INV_X1    g250(.A(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT88), .A3(G116), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n297), .A2(G122), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G107), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n202), .A3(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n433), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n196), .A2(G143), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n216), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n447), .A2(new_n449), .A3(KEYINPUT90), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT90), .B1(new_n447), .B2(new_n449), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n434), .B(new_n444), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n440), .B(KEYINPUT14), .ZN(new_n453));
  INV_X1    g267(.A(new_n439), .ZN(new_n454));
  OAI21_X1  g268(.A(G107), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n433), .B(new_n216), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n443), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n358), .A2(G217), .A3(new_n259), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n452), .B2(new_n457), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n272), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(G478), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  OAI221_X1 g280(.A(new_n272), .B1(KEYINPUT15), .B2(new_n466), .C1(new_n461), .C2(new_n462), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n259), .A2(G952), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n467), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n432), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n280), .A2(new_n356), .A3(new_n362), .A4(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n216), .A2(G137), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n219), .A2(G134), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n227), .A2(new_n197), .A3(new_n193), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT65), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n244), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n221), .A2(new_n214), .A3(new_n222), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(new_n223), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n227), .A4(new_n483), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT30), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n493), .A3(new_n484), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n309), .A2(new_n307), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n486), .A2(new_n490), .A3(new_n489), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n378), .A2(G210), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G101), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n489), .A2(new_n484), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n496), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n496), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n499), .A2(new_n509), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n505), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n507), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n491), .A2(new_n496), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n509), .B1(new_n517), .B2(new_n499), .ZN(new_n518));
  INV_X1    g332(.A(new_n511), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n506), .A2(new_n508), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G472), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n498), .B1(new_n492), .B2(new_n494), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n499), .A2(new_n529), .A3(new_n505), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n499), .A2(new_n505), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT67), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT31), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n529), .B1(new_n499), .B2(new_n505), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NOR4_X1   g351(.A1(new_n528), .A2(new_n531), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n527), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n525), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n489), .A2(new_n493), .A3(new_n484), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(KEYINPUT30), .B2(new_n491), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n534), .B(new_n530), .C1(new_n543), .C2(new_n498), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n537), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n497), .A2(KEYINPUT31), .A3(new_n534), .A4(new_n530), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n526), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n540), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n524), .B1(new_n541), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT22), .B(G137), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n295), .B2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n295), .A2(G128), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(KEYINPUT23), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT23), .B1(new_n196), .B2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n196), .A2(G119), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G110), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT68), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n557), .B2(new_n560), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n557), .A2(new_n560), .A3(new_n564), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT24), .B(G110), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n366), .B1(new_n367), .B2(new_n371), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G146), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n372), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n567), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n568), .B1(new_n575), .B2(new_n565), .ZN(new_n576));
  INV_X1    g390(.A(G110), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n558), .A2(new_n561), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n579), .A2(new_n573), .A3(new_n400), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n554), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n570), .B(new_n563), .C1(new_n373), .C2(new_n376), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n573), .A3(new_n400), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n553), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n272), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(KEYINPUT71), .A2(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n581), .A2(new_n584), .A3(new_n272), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G217), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(G234), .B2(new_n272), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n581), .A2(new_n584), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(G902), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n590), .A2(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n480), .A2(new_n550), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  OR3_X1    g411(.A1(new_n547), .A2(KEYINPUT91), .A3(G902), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT91), .B1(new_n547), .B2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(G472), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n280), .A2(new_n362), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n547), .A2(new_n548), .ZN(new_n602));
  INV_X1    g416(.A(new_n595), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n353), .A2(new_n330), .A3(new_n354), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n354), .B1(new_n353), .B2(new_n330), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n281), .B(new_n476), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n466), .A2(new_n272), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n463), .B2(G478), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n461), .B2(new_n462), .ZN(new_n611));
  INV_X1    g425(.A(new_n462), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n460), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n610), .B1(new_n615), .B2(G478), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n432), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n600), .A2(new_n601), .A3(new_n604), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND2_X1  g435(.A1(new_n539), .A2(new_n540), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n280), .A2(new_n622), .A3(new_n595), .A4(new_n362), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n539), .A2(new_n272), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(KEYINPUT91), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n623), .B1(new_n598), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT92), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n428), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n429), .A2(new_n424), .A3(new_n430), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n414), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n628), .A3(new_n414), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n465), .A2(new_n467), .B1(G475), .B2(new_n412), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n632), .A2(new_n476), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n635), .A2(KEYINPUT93), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n281), .B1(new_n605), .B2(new_n606), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n635), .B2(KEYINPUT93), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n627), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  AOI21_X1  g455(.A(new_n602), .B1(new_n626), .B2(new_n598), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n582), .A2(new_n583), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n554), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n590), .A2(new_n592), .B1(new_n594), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n479), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT37), .B(G110), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT94), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n648), .B(new_n650), .ZN(G12));
  INV_X1    g465(.A(new_n646), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n280), .A2(new_n362), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT95), .B(G900), .Z(new_n654));
  AOI21_X1  g468(.A(new_n471), .B1(new_n473), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n633), .A2(new_n632), .A3(new_n634), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n550), .A2(new_n653), .A3(new_n356), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT96), .B(G128), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G30));
  NAND2_X1  g474(.A1(new_n349), .A2(new_n355), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n661), .B(new_n662), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n405), .A2(new_n425), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT20), .ZN(new_n665));
  INV_X1    g479(.A(new_n424), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .A4(new_n427), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n630), .B2(new_n414), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n668), .A2(new_n413), .B1(new_n465), .B2(new_n467), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n281), .A2(new_n663), .A3(new_n646), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n655), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n601), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n539), .A2(new_n525), .A3(new_n540), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT32), .B1(new_n547), .B2(new_n548), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n544), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n505), .B1(new_n517), .B2(new_n499), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n272), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G472), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n670), .A2(new_n673), .A3(new_n674), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NOR2_X1   g498(.A1(new_n617), .A2(new_n655), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n550), .A2(new_n653), .A3(new_n356), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  INV_X1    g501(.A(new_n360), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n265), .A2(new_n228), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n249), .B1(new_n248), .B2(new_n254), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n261), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n233), .A2(new_n255), .A3(new_n267), .ZN(new_n692));
  AOI21_X1  g506(.A(G902), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n688), .B1(new_n693), .B2(new_n270), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n693), .B2(KEYINPUT98), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n595), .B(new_n694), .C1(new_n695), .C2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n699), .A2(new_n607), .A3(new_n617), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n550), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT41), .B(G113), .Z(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT99), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n701), .B(new_n703), .ZN(G15));
  INV_X1    g518(.A(new_n699), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n550), .A2(new_n636), .A3(new_n638), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT100), .B(G116), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G18));
  NOR3_X1   g522(.A1(new_n646), .A2(new_n432), .A3(new_n477), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n279), .A2(new_n360), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n270), .B1(new_n696), .B2(new_n697), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n693), .A2(KEYINPUT98), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n709), .A2(new_n713), .A3(new_n356), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT101), .B1(new_n550), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n624), .B1(new_n516), .B2(new_n522), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n675), .B2(new_n676), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n709), .A2(new_n713), .A3(new_n356), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n295), .ZN(G21));
  OAI21_X1  g536(.A(G472), .B1(new_n547), .B2(G902), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n506), .B1(new_n518), .B2(new_n519), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(new_n535), .B2(new_n538), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n540), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n723), .A2(new_n726), .A3(new_n595), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n661), .A2(new_n281), .A3(new_n669), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n476), .B(new_n694), .C1(new_n695), .C2(new_n698), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  AND2_X1   g546(.A1(new_n723), .A2(new_n726), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n694), .B1(new_n695), .B2(new_n698), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n637), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n652), .A3(new_n685), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  AOI21_X1  g551(.A(new_n716), .B1(new_n677), .B2(KEYINPUT103), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n675), .A2(new_n676), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n603), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n349), .A2(new_n281), .A3(new_n355), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT102), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n349), .A2(new_n744), .A3(new_n281), .A4(new_n355), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n275), .A2(G469), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n688), .B1(new_n746), .B2(new_n279), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n685), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n550), .A3(new_n595), .A4(new_n685), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n741), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n214), .ZN(G33));
  NAND4_X1  g567(.A1(new_n748), .A2(new_n550), .A3(new_n595), .A4(new_n657), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(new_n616), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n616), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n757), .A2(KEYINPUT43), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n432), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n432), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n616), .A3(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n760), .A2(new_n761), .B1(KEYINPUT43), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n652), .ZN(new_n767));
  INV_X1    g581(.A(new_n642), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n743), .A2(new_n745), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n768), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n273), .B2(new_n274), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n262), .A2(KEYINPUT45), .A3(new_n268), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(G469), .ZN(new_n778));
  NAND2_X1  g592(.A1(G469), .A2(G902), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT46), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n270), .B2(new_n693), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n779), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n688), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n671), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n771), .A2(new_n773), .A3(new_n774), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  XNOR2_X1  g600(.A(new_n783), .B(KEYINPUT47), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n717), .A2(new_n773), .A3(new_n603), .A4(new_n685), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NOR2_X1   g604(.A1(G952), .A2(G953), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT118), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n766), .A2(new_n471), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n727), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n794), .A2(KEYINPUT113), .A3(new_n772), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n794), .B2(new_n772), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n279), .B1(new_n695), .B2(new_n698), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n362), .B1(new_n797), .B2(KEYINPUT115), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n795), .B(new_n796), .C1(new_n787), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n772), .A2(new_n734), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n652), .A2(new_n793), .A3(new_n733), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n682), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n803), .A3(new_n595), .A4(new_n471), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n432), .A3(new_n616), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n663), .A2(new_n281), .A3(new_n734), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n766), .A3(new_n471), .A4(new_n727), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n808), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n793), .A2(new_n735), .A3(new_n727), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n816), .B(new_n468), .C1(new_n617), .C2(new_n806), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n793), .A2(new_n741), .A3(new_n803), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n818), .A2(KEYINPUT48), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(KEYINPUT48), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n812), .A2(KEYINPUT116), .A3(new_n813), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT116), .B1(new_n812), .B2(new_n813), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n808), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n808), .B(KEYINPUT117), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n800), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n795), .B(new_n796), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n815), .B(new_n821), .C1(new_n832), .C2(KEYINPUT51), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n747), .A2(new_n646), .A3(new_n656), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n728), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n682), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n658), .A2(new_n686), .A3(new_n837), .A4(new_n736), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n550), .A2(new_n700), .B1(new_n727), .B2(new_n730), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n706), .C1(new_n715), .C2(new_n720), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n413), .A2(new_n465), .A3(new_n467), .A4(new_n656), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n632), .A3(new_n633), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT108), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n632), .A3(KEYINPUT108), .A4(new_n633), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n773), .A2(new_n848), .A3(new_n550), .A4(new_n653), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n733), .A2(new_n652), .A3(new_n685), .ZN(new_n850));
  INV_X1    g664(.A(new_n748), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n849), .B(new_n754), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n752), .A2(new_n842), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n465), .A2(new_n467), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n761), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n607), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n627), .A2(new_n856), .B1(new_n642), .B2(new_n647), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT107), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n596), .A4(new_n619), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n600), .A2(new_n601), .A3(new_n856), .A4(new_n604), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n648), .A2(new_n619), .A3(new_n860), .A4(new_n596), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT107), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n840), .A2(new_n853), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n834), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n834), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n838), .A2(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n658), .A2(new_n736), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n873), .A2(KEYINPUT109), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(KEYINPUT109), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n686), .A3(new_n837), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n876), .B2(KEYINPUT52), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n842), .B(KEYINPUT111), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n752), .A2(new_n852), .A3(new_n865), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n863), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n864), .A2(new_n834), .A3(new_n865), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n880), .B(new_n871), .C1(new_n882), .C2(new_n866), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT112), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n853), .A2(new_n863), .A3(new_n865), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n885), .A2(new_n877), .B1(new_n864), .B2(KEYINPUT53), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n881), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n792), .B1(new_n833), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT106), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n595), .A2(new_n362), .A3(new_n281), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n663), .A2(new_n765), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n805), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n891), .B2(new_n895), .ZN(G75));
  AOI21_X1  g710(.A(new_n272), .B1(new_n869), .B2(new_n880), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT120), .A3(new_n348), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n880), .B1(new_n882), .B2(new_n866), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(G902), .A3(new_n348), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n342), .B(KEYINPUT119), .Z(new_n903));
  XOR2_X1   g717(.A(new_n344), .B(KEYINPUT55), .Z(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n898), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n259), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n900), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n905), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n907), .A2(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n883), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n899), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n779), .B(KEYINPUT57), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n691), .A2(new_n692), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n921));
  INV_X1    g735(.A(new_n778), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n897), .B2(new_n922), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n921), .A2(new_n899), .A3(G902), .A4(new_n922), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n908), .B1(new_n920), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  INV_X1    g741(.A(new_n426), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n908), .ZN(G60));
  INV_X1    g745(.A(new_n615), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n608), .B(KEYINPUT59), .Z(new_n933));
  NAND4_X1  g747(.A1(new_n915), .A2(new_n932), .A3(new_n916), .A4(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n908), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n888), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n645), .B(KEYINPUT124), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n899), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n899), .A2(new_n941), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n935), .B(new_n943), .C1(new_n944), .C2(new_n593), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G66));
  INV_X1    g761(.A(G224), .ZN(new_n948));
  OAI21_X1  g762(.A(G953), .B1(new_n474), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n863), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n842), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n903), .B1(G898), .B2(new_n259), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  AND3_X1   g768(.A1(new_n874), .A2(new_n686), .A3(new_n875), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n683), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n772), .B(new_n672), .C1(new_n617), .C2(new_n855), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n550), .A3(new_n595), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n785), .A2(new_n789), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n259), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n421), .B(KEYINPUT125), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n495), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n784), .A2(new_n356), .A3(new_n669), .A4(new_n741), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n789), .A2(new_n754), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n752), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n785), .A2(new_n968), .A3(new_n969), .A4(new_n955), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(G953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n972));
  AOI22_X1  g786(.A1(new_n963), .A2(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  INV_X1    g791(.A(new_n951), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n962), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n505), .A3(new_n500), .ZN(new_n980));
  INV_X1    g794(.A(new_n977), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n507), .B2(new_n544), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT126), .Z(new_n983));
  NAND2_X1  g797(.A1(new_n886), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n977), .B1(new_n970), .B2(new_n978), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n500), .A2(new_n505), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n908), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n980), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n980), .A2(new_n984), .A3(new_n990), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(G57));
endmodule


