//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  INV_X1    g0004(.A(G58), .ZN(new_n205));
  INV_X1    g0005(.A(G232), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(G238), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n209), .B1(G68), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G97), .A2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  NAND3_X1  g0020(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n223));
  OAI21_X1  g0023(.A(G20), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n203), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  AND2_X1   g0029(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n230));
  NOR4_X1   g0030(.A1(new_n220), .A2(new_n226), .A3(new_n229), .A4(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT67), .B(G250), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G257), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n206), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT16), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT7), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n253), .A4(new_n254), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n205), .A2(new_n249), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G58), .A2(G68), .ZN(new_n261));
  OAI21_X1  g0061(.A(G20), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G159), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n248), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT75), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT64), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n270), .A2(new_n221), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n257), .A2(new_n258), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n265), .B1(new_n273), .B2(G68), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(KEYINPUT16), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT75), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n276), .B(new_n248), .C1(new_n259), .C2(new_n265), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n267), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n272), .B1(G1), .B2(new_n253), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n222), .A2(new_n223), .B1(new_n251), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  AND2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n291), .B1(G223), .B2(G1698), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G87), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n281), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(G1), .B(G13), .C1(new_n251), .C2(new_n288), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n297), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n300), .B1(new_n302), .B2(new_n206), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n296), .A2(new_n303), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(G200), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n278), .A2(new_n287), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT76), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n278), .A2(new_n310), .A3(new_n307), .A4(new_n287), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n292), .A2(new_n293), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT7), .B1(new_n313), .B2(new_n253), .ZN(new_n314));
  INV_X1    g0114(.A(new_n258), .ZN(new_n315));
  OAI21_X1  g0115(.A(G68), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n265), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n276), .B1(new_n318), .B2(new_n248), .ZN(new_n319));
  INV_X1    g0119(.A(new_n277), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n286), .B1(new_n321), .B2(new_n275), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(KEYINPUT77), .A3(new_n323), .A4(new_n307), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n278), .A2(new_n323), .A3(new_n307), .A4(new_n287), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT77), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(KEYINPUT17), .A2(new_n312), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n252), .A2(new_n254), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G222), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G223), .A2(G1698), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n270), .A2(new_n221), .B1(G33), .B2(G41), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n335), .C1(G77), .C2(new_n330), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(new_n300), .C1(new_n290), .C2(new_n302), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G200), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT69), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n304), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n270), .A2(new_n221), .A3(new_n271), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n251), .A2(G20), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n279), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G150), .ZN(new_n346));
  INV_X1    g0146(.A(new_n263), .ZN(new_n347));
  NOR3_X1   g0147(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n346), .A2(new_n347), .B1(new_n348), .B2(new_n253), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n285), .A2(G50), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  INV_X1    g0152(.A(G50), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n282), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n351), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT9), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n341), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT10), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT10), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n341), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n278), .A2(new_n287), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n306), .A2(G169), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n306), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT18), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n337), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n357), .B(new_n372), .C1(G179), .C2(new_n337), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n329), .A2(new_n363), .A3(new_n370), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n290), .A2(new_n331), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n330), .B(new_n375), .C1(G232), .C2(new_n331), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT70), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(G33), .A3(G97), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n289), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n300), .B1(new_n302), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT13), .B1(new_n382), .B2(new_n386), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(KEYINPUT71), .A3(new_n389), .ZN(new_n390));
  OR4_X1    g0190(.A1(KEYINPUT71), .A2(new_n382), .A3(KEYINPUT13), .A4(new_n386), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(G169), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT73), .B(KEYINPUT14), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n390), .A2(new_n391), .A3(G169), .A4(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(G179), .A3(new_n389), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n394), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n343), .A2(G77), .B1(G20), .B2(new_n249), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n353), .B2(new_n347), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n403), .A2(new_n342), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n404), .A2(KEYINPUT11), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(KEYINPUT11), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n283), .A2(new_n249), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT12), .ZN(new_n408));
  INV_X1    g0208(.A(new_n285), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n405), .A2(new_n406), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n388), .A2(G190), .A3(new_n389), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n411), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n390), .A2(new_n391), .A3(G200), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n280), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT15), .B(G87), .Z(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n344), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n342), .B1(new_n409), .B2(G77), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G77), .B2(new_n282), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n330), .B1(new_n206), .B2(G1698), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n210), .A2(new_n331), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n335), .B1(G107), .B2(new_n330), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n302), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n299), .B1(new_n428), .B2(G244), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n366), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n424), .B(new_n432), .C1(G169), .C2(new_n431), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n412), .A2(new_n418), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n424), .B1(G190), .B2(new_n431), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n431), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n374), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT24), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n253), .B(G87), .C1(new_n292), .C2(new_n293), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT22), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n330), .A2(KEYINPUT22), .A3(new_n253), .A4(G87), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  INV_X1    g0246(.A(G107), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(G20), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT85), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n450), .A2(new_n446), .A3(new_n447), .A4(G20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n453), .A2(G20), .B1(new_n446), .B2(new_n447), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n440), .B1(new_n445), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n449), .B2(new_n451), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(KEYINPUT24), .A3(new_n443), .A4(new_n444), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n342), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT86), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT25), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n464));
  NOR4_X1   g0264(.A1(new_n463), .A2(new_n282), .A3(G107), .A4(new_n464), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n461), .B(new_n462), .C1(new_n283), .C2(new_n447), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n251), .B2(G1), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(new_n270), .A3(new_n221), .A4(new_n271), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n281), .A2(KEYINPUT78), .A3(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n282), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI211_X1 g0272(.A(new_n465), .B(new_n466), .C1(G107), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n460), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n330), .B1(G257), .B2(new_n331), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G250), .A2(G1698), .ZN(new_n476));
  INV_X1    g0276(.A(G294), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n475), .A2(new_n476), .B1(new_n251), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n335), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(new_n301), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n484), .A2(new_n298), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n479), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n371), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n479), .A2(new_n366), .A3(new_n486), .A4(new_n487), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n474), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT87), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n474), .A2(new_n489), .A3(new_n493), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n488), .A2(new_n304), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n474), .ZN(new_n497));
  INV_X1    g0297(.A(new_n488), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n436), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n472), .A2(new_n420), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n378), .A2(new_n380), .A3(KEYINPUT19), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n253), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n214), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n330), .A2(new_n253), .A3(G68), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT19), .B1(new_n343), .B2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n342), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n420), .A2(new_n282), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n502), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n504), .B2(new_n506), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n272), .B1(new_n516), .B2(new_n508), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n517), .A2(KEYINPUT81), .A3(new_n513), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n501), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n481), .A2(new_n298), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n215), .B1(new_n480), .B2(G1), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n301), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n208), .A2(G1698), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n523), .B1(G238), .B2(G1698), .C1(new_n292), .C2(new_n293), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G179), .B(new_n522), .C1(new_n526), .C2(new_n289), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n289), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  INV_X1    g0328(.A(new_n522), .ZN(new_n529));
  OAI21_X1  g0329(.A(G169), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT80), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n527), .B2(new_n530), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n472), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n214), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT81), .B1(new_n517), .B2(new_n513), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n503), .A2(new_n253), .B1(new_n214), .B2(new_n505), .ZN(new_n538));
  INV_X1    g0338(.A(new_n508), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(new_n509), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n502), .B(new_n514), .C1(new_n540), .C2(new_n272), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n536), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n528), .A2(new_n529), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n304), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G200), .B2(new_n543), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n519), .A2(new_n534), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(new_n331), .C1(new_n292), .C2(new_n293), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT79), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT4), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n330), .A2(G244), .A3(new_n331), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G283), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n330), .A2(G250), .A3(G1698), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n335), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n484), .A2(G257), .A3(new_n301), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n487), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n273), .A2(G107), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  AND2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n505), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n447), .A2(KEYINPUT6), .A3(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n272), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n535), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n282), .A2(G97), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n557), .B1(new_n555), .B2(new_n335), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(G190), .A3(new_n487), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n560), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n559), .A2(new_n371), .ZN(new_n576));
  INV_X1    g0376(.A(new_n566), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n577), .A2(new_n253), .B1(new_n207), .B2(new_n347), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n447), .B1(new_n257), .B2(new_n258), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n342), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n570), .ZN(new_n581));
  INV_X1    g0381(.A(new_n571), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n573), .A2(new_n366), .A3(new_n487), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n546), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n553), .B(new_n253), .C1(G33), .C2(new_n569), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G20), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n342), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT20), .ZN(new_n592));
  INV_X1    g0392(.A(new_n471), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n272), .A2(new_n593), .A3(G116), .A4(new_n468), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT20), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n342), .A2(new_n595), .A3(new_n588), .A4(new_n590), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n282), .A2(G116), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n592), .A2(new_n594), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n597), .B1(new_n472), .B2(G116), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(KEYINPUT82), .A3(new_n592), .A4(new_n596), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G303), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n313), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n331), .A2(G257), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G264), .A2(G1698), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n292), .C2(new_n293), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(new_n335), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n484), .A2(G270), .A3(new_n301), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n487), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G169), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n604), .A2(new_n618), .A3(new_n614), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n613), .A2(new_n617), .B1(new_n366), .B2(new_n612), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n604), .A2(new_n621), .A3(KEYINPUT83), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT83), .B1(new_n604), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n612), .A2(new_n304), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(G200), .B2(new_n612), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n601), .A3(new_n603), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n620), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n439), .A2(new_n500), .A3(new_n587), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT88), .ZN(G372));
  INV_X1    g0430(.A(new_n418), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n412), .B2(new_n433), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n369), .B1(new_n632), .B2(new_n329), .ZN(new_n633));
  INV_X1    g0433(.A(new_n363), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n373), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(KEYINPUT90), .B(new_n373), .C1(new_n633), .C2(new_n634), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n439), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n546), .A2(KEYINPUT26), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT89), .ZN(new_n643));
  INV_X1    g0443(.A(new_n536), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n644), .B(new_n545), .C1(new_n515), .C2(new_n518), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n537), .A2(new_n541), .B1(new_n472), .B2(new_n420), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n527), .A2(new_n530), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n641), .B(new_n645), .C1(new_n646), .C2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n546), .A2(new_n652), .A3(KEYINPUT26), .A4(new_n641), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n643), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n519), .A2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n604), .A2(new_n621), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n620), .A2(new_n491), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n586), .A2(new_n499), .A3(new_n645), .A4(new_n655), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n639), .B1(new_n640), .B2(new_n660), .ZN(G369));
  NAND2_X1  g0461(.A1(new_n620), .A2(new_n656), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n253), .A2(G13), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .A3(G1), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT27), .B1(new_n663), .B2(G1), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n604), .A2(new_n668), .ZN(new_n669));
  MUX2_X1   g0469(.A(new_n662), .B(new_n628), .S(new_n669), .Z(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n474), .A2(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n500), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n668), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n491), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n491), .A2(new_n668), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n668), .B1(new_n620), .B2(new_n624), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n500), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n227), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n506), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n225), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(new_n655), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n546), .A2(new_n650), .A3(new_n641), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n495), .A2(new_n620), .A3(new_n624), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n658), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n693), .A2(KEYINPUT91), .A3(new_n675), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT91), .B1(new_n693), .B2(new_n675), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT29), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n660), .B2(new_n668), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n488), .A2(new_n612), .ZN(new_n700));
  INV_X1    g0500(.A(new_n527), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n573), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n498), .A2(new_n543), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n366), .A3(new_n559), .A4(new_n612), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n700), .A2(KEYINPUT30), .A3(new_n701), .A4(new_n573), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n668), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n495), .A2(new_n546), .A3(new_n586), .A4(new_n499), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n620), .A2(new_n624), .A3(new_n627), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n668), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n699), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n688), .B1(new_n719), .B2(G1), .ZN(G364));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n670), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n270), .A2(new_n221), .B1(G20), .B2(new_n371), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n366), .A2(new_n436), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n253), .A2(G190), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n249), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n436), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n447), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G159), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT32), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n253), .A2(new_n304), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n731), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G87), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n727), .A2(new_n739), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n353), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n253), .B1(new_n734), .B2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n366), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n728), .A2(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n330), .B1(new_n745), .B2(new_n569), .C1(new_n207), .C2(new_n747), .ZN(new_n748));
  OR4_X1    g0548(.A1(new_n733), .A2(new_n738), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n739), .A2(new_n746), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n730), .B(new_n749), .C1(G58), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n729), .ZN(new_n753));
  INV_X1    g0553(.A(G317), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n736), .A2(G329), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n732), .ZN(new_n760));
  INV_X1    g0560(.A(new_n743), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(G326), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n741), .A2(G303), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n330), .B1(new_n751), .B2(G322), .ZN(new_n764));
  INV_X1    g0564(.A(new_n745), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G294), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n747), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G311), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n726), .B1(new_n752), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n682), .A2(new_n330), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G45), .B2(new_n225), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n480), .B2(new_n243), .ZN(new_n774));
  INV_X1    g0574(.A(G355), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n330), .A2(new_n227), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(G116), .B2(new_n227), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n726), .A2(new_n723), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n663), .B(KEYINPUT93), .Z(new_n780));
  AOI21_X1  g0580(.A(new_n281), .B1(new_n780), .B2(G45), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n683), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n725), .A2(new_n770), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n672), .A2(KEYINPUT92), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n670), .A2(G330), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n784), .B1(new_n787), .B2(new_n783), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n424), .A2(new_n668), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n437), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n433), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n433), .A2(new_n668), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n660), .B2(new_n668), .ZN(new_n795));
  INV_X1    g0595(.A(new_n794), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n675), .B(new_n796), .C1(new_n654), .C2(new_n659), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(new_n717), .ZN(new_n799));
  INV_X1    g0599(.A(new_n783), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n794), .A2(new_n721), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n726), .A2(new_n721), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n207), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G143), .A2(new_n751), .B1(new_n768), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n806), .B2(new_n743), .C1(new_n346), .C2(new_n729), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT34), .Z(new_n808));
  NOR2_X1   g0608(.A1(new_n732), .A2(new_n249), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G50), .B2(new_n741), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n313), .B1(new_n765), .B2(G58), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n735), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n729), .A2(new_n759), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n313), .B1(new_n740), .B2(new_n447), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT95), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n751), .A2(G294), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n743), .A2(new_n605), .B1(new_n745), .B2(new_n569), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G116), .B2(new_n768), .ZN(new_n820));
  INV_X1    g0620(.A(new_n732), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G87), .A2(new_n821), .B1(new_n736), .B2(G311), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n808), .A2(new_n814), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n726), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n802), .A2(new_n783), .A3(new_n804), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n801), .A2(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n412), .A2(new_n668), .ZN(new_n828));
  INV_X1    g0628(.A(new_n666), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n275), .A2(new_n266), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n287), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(new_n328), .C2(new_n369), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT97), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n368), .B(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n364), .A2(new_n829), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n312), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n367), .A2(new_n829), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n309), .A2(new_n311), .B1(new_n838), .B2(new_n831), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n834), .A2(new_n837), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT38), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n832), .A2(KEYINPUT38), .A3(new_n840), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(KEYINPUT39), .A3(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n832), .A2(KEYINPUT38), .A3(new_n840), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n325), .B(KEYINPUT77), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n323), .B1(new_n309), .B2(new_n311), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT100), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n312), .A2(KEYINPUT17), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n324), .A2(new_n327), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n848), .A2(new_n852), .A3(new_n370), .ZN(new_n853));
  INV_X1    g0653(.A(new_n836), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n368), .A2(new_n836), .A3(new_n308), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT99), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT37), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n368), .B(KEYINPUT97), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n861), .A2(new_n835), .A3(new_n312), .A4(new_n836), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n845), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n828), .B(new_n844), .C1(new_n866), .C2(KEYINPUT39), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n412), .B(new_n418), .C1(new_n416), .C2(new_n675), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n401), .A2(new_n411), .A3(new_n668), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n797), .B2(new_n793), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n842), .A2(new_n843), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n872), .A2(new_n873), .B1(new_n369), .B2(new_n666), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n696), .A2(new_n698), .A3(new_n439), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n639), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n875), .B(new_n877), .Z(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n715), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n714), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n794), .B1(new_n868), .B2(new_n869), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT40), .B1(new_n866), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n709), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n628), .A2(new_n500), .A3(new_n587), .A4(new_n675), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(KEYINPUT31), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n715), .B(KEYINPUT101), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n883), .B(new_n888), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n873), .B2(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n439), .A3(new_n882), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n883), .B1(new_n891), .B2(new_n892), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT102), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n853), .A2(new_n854), .B1(new_n860), .B2(new_n862), .ZN(new_n900));
  INV_X1    g0700(.A(new_n865), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n843), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n886), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n845), .A2(new_n841), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n893), .B1(new_n904), .B2(new_n886), .ZN(new_n905));
  OAI21_X1  g0705(.A(G330), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(G330), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n714), .B2(new_n881), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n439), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n897), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n878), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n281), .B2(new_n780), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT35), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n224), .B1(new_n577), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(G116), .C1(new_n914), .C2(new_n577), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT36), .ZN(new_n917));
  OAI21_X1  g0717(.A(G77), .B1(new_n205), .B2(new_n249), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n918), .A2(new_n225), .B1(G50), .B2(new_n249), .ZN(new_n919));
  INV_X1    g0719(.A(G13), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(G1), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n913), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT103), .Z(G367));
  XNOR2_X1  g0723(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n500), .A2(new_n679), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n575), .A2(new_n585), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n583), .B2(new_n668), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT42), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n585), .B1(new_n928), .B2(new_n495), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n675), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n655), .A2(new_n645), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n542), .A2(new_n675), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n655), .ZN(new_n938));
  MUX2_X1   g0738(.A(new_n937), .B(new_n934), .S(new_n938), .Z(new_n939));
  INV_X1    g0739(.A(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n933), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n930), .A2(new_n940), .A3(new_n939), .A4(new_n932), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n924), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(new_n924), .A3(new_n944), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n641), .A2(new_n668), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n677), .B1(new_n928), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n948), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n925), .B1(new_n676), .B2(new_n679), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n671), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n677), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n718), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n928), .A2(new_n949), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n680), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT44), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n680), .A2(new_n958), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n957), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n719), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n683), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n782), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n939), .A2(new_n723), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n761), .A2(G143), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n821), .A2(G77), .ZN(new_n972));
  INV_X1    g0772(.A(G159), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n729), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n750), .A2(new_n346), .B1(new_n745), .B2(new_n249), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n974), .A2(new_n313), .A3(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n740), .A2(new_n205), .B1(new_n735), .B2(new_n806), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT107), .Z(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(new_n353), .C2(new_n747), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n741), .A2(G116), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT46), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n750), .A2(new_n605), .B1(new_n735), .B2(new_n754), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G97), .B2(new_n821), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G294), .A2(new_n753), .B1(new_n768), .B2(G283), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n330), .B1(new_n765), .B2(G107), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n981), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(G311), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n743), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n979), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n726), .ZN(new_n991));
  INV_X1    g0791(.A(new_n771), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n235), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n778), .B1(new_n227), .B2(new_n421), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n991), .B(new_n783), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT108), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n952), .A2(new_n969), .B1(new_n970), .B2(new_n996), .ZN(G387));
  NAND2_X1  g0797(.A1(new_n955), .A2(new_n782), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT109), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n676), .A2(new_n724), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n421), .A2(new_n745), .B1(new_n973), .B2(new_n743), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n740), .A2(new_n207), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G97), .B2(new_n821), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1003), .B(new_n330), .C1(new_n346), .C2(new_n735), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT111), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1001), .B(new_n1005), .C1(G50), .C2(new_n751), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n249), .B2(new_n747), .C1(new_n279), .C2(new_n729), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G311), .A2(new_n753), .B1(new_n751), .B2(G317), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(KEYINPUT112), .B(G322), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n761), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(new_n605), .C2(new_n747), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT48), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n759), .B2(new_n745), .C1(new_n477), .C2(new_n740), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT49), .Z(new_n1014));
  AOI21_X1  g0814(.A(new_n330), .B1(new_n736), .B2(G326), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n589), .B2(new_n732), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1007), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n726), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n239), .A2(G45), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT110), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n279), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g0822(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n685), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1020), .A2(new_n771), .A3(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(G107), .B2(new_n227), .C1(new_n685), .C2(new_n776), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n778), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1000), .A2(new_n1018), .A3(new_n783), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n719), .A2(new_n955), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n683), .B1(new_n956), .B2(new_n718), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n999), .B(new_n1028), .C1(new_n1029), .C2(new_n1030), .ZN(G393));
  INV_X1    g0831(.A(KEYINPUT113), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n964), .B(new_n961), .C1(new_n1032), .C2(new_n677), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n677), .A2(new_n1032), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1033), .B(new_n1034), .Z(new_n1035));
  OAI211_X1 g0835(.A(new_n683), .B(new_n966), .C1(new_n1035), .C2(new_n957), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n313), .B1(new_n736), .B2(G143), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n249), .B2(new_n740), .C1(new_n214), .C2(new_n732), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT115), .Z(new_n1039));
  OAI22_X1  g0839(.A1(new_n743), .A2(new_n346), .B1(new_n750), .B2(new_n973), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT114), .Z(new_n1041));
  AOI22_X1  g0841(.A1(new_n1041), .A2(KEYINPUT51), .B1(G77), .B2(new_n765), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(KEYINPUT51), .B2(new_n1041), .C1(new_n279), .C2(new_n747), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1039), .B(new_n1043), .C1(G50), .C2(new_n753), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n743), .A2(new_n754), .B1(new_n750), .B2(new_n987), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n741), .A2(G283), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n745), .A2(new_n589), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1048), .B(new_n733), .C1(G303), .C2(new_n753), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n330), .B1(new_n736), .B2(new_n1009), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G294), .B2(new_n768), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n726), .B1(new_n1044), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n928), .A2(new_n723), .A3(new_n949), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n778), .B1(new_n569), .B2(new_n227), .C1(new_n246), .C2(new_n992), .ZN(new_n1055));
  AND4_X1   g0855(.A1(new_n783), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1035), .B2(new_n782), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1036), .A2(new_n1057), .ZN(G390));
  NAND2_X1  g0858(.A1(new_n908), .A2(new_n883), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n693), .A2(new_n675), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT91), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n693), .A2(KEYINPUT91), .A3(new_n675), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n793), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(new_n791), .A3(new_n870), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n828), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1065), .A2(new_n902), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT39), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n902), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n797), .A2(new_n793), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n870), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1069), .A2(new_n844), .B1(new_n1071), .B2(new_n1066), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1059), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1069), .A2(new_n844), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1066), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1065), .A2(new_n902), .A3(new_n1066), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n716), .A2(G330), .A3(new_n796), .A4(new_n870), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1073), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n694), .A2(new_n695), .A3(new_n792), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n791), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n870), .B1(new_n908), .B2(new_n796), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n715), .ZN(new_n1086));
  OAI211_X1 g0886(.A(G330), .B(new_n796), .C1(new_n891), .C2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(new_n871), .B1(new_n908), .B2(new_n883), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1070), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1084), .A2(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n876), .A2(new_n639), .A3(new_n909), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1081), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1073), .A2(new_n1080), .A3(new_n1092), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n683), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1074), .A2(new_n721), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n753), .A2(G137), .B1(new_n765), .B2(G159), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n747), .B2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT116), .Z(new_n1102));
  NOR2_X1   g0902(.A1(new_n740), .A2(new_n346), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n313), .B1(new_n821), .B2(G50), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G128), .B2(new_n761), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n735), .C1(new_n813), .C2(new_n750), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT117), .Z(new_n1110));
  OAI221_X1 g0910(.A(new_n742), .B1(new_n735), .B2(new_n477), .C1(new_n569), .C2(new_n747), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n809), .B(new_n1111), .C1(G107), .C2(new_n753), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n750), .A2(new_n589), .B1(new_n745), .B2(new_n207), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT118), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n313), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G283), .B2(new_n761), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n726), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n803), .A2(new_n279), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1097), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1081), .A2(new_n782), .B1(new_n783), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1096), .A2(new_n1120), .ZN(G378));
  NAND3_X1  g0921(.A1(new_n906), .A2(new_n867), .A3(new_n874), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n875), .A2(new_n896), .A3(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n363), .A2(new_n373), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT121), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n357), .A2(new_n829), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1122), .A2(new_n1123), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n782), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n353), .B1(new_n292), .B2(G41), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n747), .A2(new_n806), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1100), .A2(new_n740), .B1(new_n346), .B2(new_n745), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(G128), .C2(new_n751), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n1108), .B2(new_n743), .C1(new_n813), .C2(new_n729), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G41), .B1(new_n736), .B2(G124), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n251), .C1(new_n973), .C2(new_n732), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1137), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n288), .B1(new_n735), .B2(new_n759), .C1(new_n447), .C2(new_n750), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n743), .A2(new_n589), .B1(new_n745), .B2(new_n249), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1002), .B(new_n1147), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n313), .B1(new_n729), .B2(new_n569), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n420), .B2(new_n768), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n205), .C2(new_n732), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT58), .Z(new_n1155));
  OAI21_X1  g0955(.A(new_n726), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n800), .B1(new_n353), .B2(new_n803), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1133), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1156), .B(new_n1157), .C1(new_n1158), .C2(new_n722), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1136), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1092), .B1(new_n1073), .B2(new_n1080), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n876), .A2(new_n639), .A3(new_n909), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1134), .A2(new_n1135), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT57), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n683), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1158), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1122), .A2(new_n1123), .A3(new_n1133), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1094), .A2(new_n1091), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1160), .B1(new_n1165), .B2(new_n1171), .ZN(G375));
  INV_X1    g0972(.A(new_n1090), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1162), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n968), .A3(new_n1092), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n972), .B1(new_n759), .B2(new_n750), .C1(new_n421), .C2(new_n745), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n761), .A2(G294), .B1(new_n768), .B2(G107), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n589), .B2(new_n729), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT122), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT122), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n330), .B(new_n1176), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n569), .B2(new_n740), .C1(new_n605), .C2(new_n735), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT123), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n330), .B1(new_n735), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G137), .A2(new_n751), .B1(new_n821), .B2(G58), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n813), .B2(new_n743), .C1(new_n346), .C2(new_n747), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G159), .C2(new_n741), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n353), .B2(new_n745), .C1(new_n729), .C2(new_n1100), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n800), .B1(new_n1191), .B2(new_n726), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n722), .B2(new_n870), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n249), .B2(new_n803), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1090), .B2(new_n782), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1175), .A2(new_n1195), .ZN(G381));
  XOR2_X1   g0996(.A(G375), .B(KEYINPUT124), .Z(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(G378), .ZN(new_n1198));
  INV_X1    g0998(.A(G384), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n1195), .A4(new_n1175), .ZN(new_n1200));
  OR2_X1    g1000(.A1(G387), .A2(G390), .ZN(new_n1201));
  OR3_X1    g1001(.A1(new_n1201), .A2(G396), .A3(G393), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1200), .A2(new_n1202), .ZN(G407));
  INV_X1    g1003(.A(G213), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1198), .B2(new_n667), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1200), .B2(new_n1202), .ZN(G409));
  NOR2_X1   g1006(.A1(new_n1204), .A2(G343), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G378), .B(new_n1160), .C1(new_n1165), .C2(new_n1171), .ZN(new_n1208));
  INV_X1    g1008(.A(G378), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n968), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1163), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1136), .A2(new_n1159), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1209), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1207), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n684), .B1(new_n1174), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n1092), .C1(new_n1216), .C2(new_n1174), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(G384), .A3(new_n1195), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G384), .B1(new_n1218), .B2(new_n1195), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1214), .A2(new_n1215), .A3(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(G393), .B(G396), .Z(new_n1224));
  NAND2_X1  g1024(.A1(G387), .A2(G390), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G387), .A2(G390), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1224), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1201), .A2(new_n1229), .A3(new_n1225), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT61), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G2897), .B(new_n1207), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1221), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1207), .A2(G2897), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1219), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1223), .B(new_n1231), .C1(new_n1214), .C2(new_n1236), .ZN(new_n1237));
  AND2_X1   g1037(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1215), .B(new_n1238), .C1(new_n1214), .C2(new_n1222), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1207), .ZN(new_n1242));
  AND4_X1   g1042(.A1(KEYINPUT63), .A2(new_n1241), .A3(new_n1242), .A4(new_n1222), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT63), .B1(new_n1214), .B2(new_n1222), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1236), .B2(new_n1214), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1236), .A2(new_n1214), .A3(new_n1247), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1240), .B1(new_n1250), .B2(new_n1252), .ZN(G405));
  NAND2_X1  g1053(.A1(G375), .A2(new_n1209), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1208), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(new_n1222), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(new_n1251), .ZN(G402));
endmodule


