//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G134), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT66), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT68), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n197));
  AOI21_X1  g011(.A(G137), .B1(new_n190), .B2(new_n192), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n197), .B(G131), .C1(new_n198), .C2(new_n188), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n191), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n189), .A2(KEYINPUT66), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n201), .B(new_n187), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n201), .B1(G134), .B2(new_n187), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n190), .A2(new_n192), .A3(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(G134), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G137), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n195), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n200), .A2(KEYINPUT73), .A3(new_n213), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT64), .A2(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT64), .A2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(G146), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n220), .A2(G128), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  INV_X1    g039(.A(new_n221), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n223), .ZN(new_n227));
  AOI21_X1  g041(.A(G146), .B1(new_n218), .B2(new_n219), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n222), .A2(G143), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n224), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n216), .A2(new_n217), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n228), .B2(new_n229), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT65), .B(new_n235), .C1(new_n228), .C2(new_n229), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n220), .A2(new_n223), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n238), .A2(new_n239), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n209), .A2(new_n212), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n205), .B1(new_n198), .B2(new_n201), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n244), .A2(KEYINPUT72), .A3(new_n213), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT72), .B1(new_n244), .B2(new_n213), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G116), .B(G119), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT2), .A2(G113), .ZN(new_n250));
  AND3_X1   g064(.A1(KEYINPUT71), .A2(KEYINPUT2), .A3(G113), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT71), .B1(KEYINPUT2), .B2(G113), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n248), .B(new_n250), .C1(new_n252), .C2(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n232), .A2(new_n247), .A3(new_n257), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT74), .B(KEYINPUT27), .Z(new_n259));
  INV_X1    g073(.A(G237), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n259), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n263), .B(new_n264), .Z(new_n265));
  NAND2_X1  g079(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(KEYINPUT75), .A3(new_n265), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n232), .A2(new_n247), .A3(KEYINPUT30), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n200), .A2(new_n213), .A3(new_n231), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n200), .A2(new_n273), .A3(new_n231), .A4(new_n213), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n244), .A2(new_n213), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n241), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n279), .A3(new_n256), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n268), .A2(new_n269), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT31), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n258), .A2(KEYINPUT28), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n232), .A2(new_n247), .A3(new_n284), .A4(new_n257), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n277), .A2(new_n256), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n265), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n268), .A2(new_n291), .A3(new_n269), .A4(new_n280), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n282), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n296), .A2(G472), .A3(G902), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n283), .A2(new_n285), .B1(new_n256), .B2(new_n277), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n292), .B1(new_n265), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n270), .A2(new_n279), .A3(new_n256), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT75), .B1(new_n258), .B2(new_n265), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n291), .B1(new_n303), .B2(new_n269), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n298), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n257), .B1(new_n232), .B2(new_n247), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n283), .B2(new_n285), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n289), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n286), .A2(new_n313), .A3(new_n265), .A4(new_n287), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n280), .A2(new_n258), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n289), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n310), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n299), .B2(new_n265), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G472), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n293), .A2(KEYINPUT77), .A3(new_n298), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n297), .A2(new_n307), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G469), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n261), .A2(G227), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G107), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G104), .ZN(new_n330));
  INV_X1    g144(.A(G104), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT85), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n330), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(G101), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n231), .A3(KEYINPUT10), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n339), .B1(new_n330), .B2(new_n332), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n338), .A2(KEYINPUT85), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n347), .A2(new_n335), .B1(G104), .B2(new_n329), .ZN(new_n348));
  OAI21_X1  g162(.A(G101), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n342), .A3(KEYINPUT4), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n351), .B(G101), .C1(new_n346), .C2(new_n348), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n241), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT86), .ZN(new_n354));
  AND2_X1   g168(.A1(KEYINPUT64), .A2(G143), .ZN(new_n355));
  NOR2_X1   g169(.A1(KEYINPUT64), .A2(G143), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n222), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n225), .B1(new_n357), .B2(KEYINPUT1), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n224), .B1(new_n240), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n344), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT86), .B(KEYINPUT10), .C1(new_n344), .C2(new_n359), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n345), .B(new_n353), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n245), .A2(new_n246), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n328), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT72), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n275), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n244), .A2(new_n213), .A3(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n342), .A2(new_n343), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n371), .B(new_n224), .C1(new_n230), .C2(new_n227), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n369), .A2(new_n370), .B1(new_n360), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT87), .B1(new_n373), .B2(KEYINPUT12), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n360), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n245), .B2(new_n246), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n367), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n364), .A2(new_n366), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n353), .A2(new_n345), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(new_n365), .C1(new_n363), .C2(new_n362), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n328), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n323), .B(new_n324), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n367), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n383), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n364), .A2(new_n366), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n380), .B2(new_n381), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n389), .B(G469), .C1(new_n391), .C2(new_n328), .ZN(new_n392));
  NAND2_X1  g206(.A1(G469), .A2(G902), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  OAI21_X1  g209(.A(G221), .B1(new_n395), .B2(G902), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G214), .B1(G237), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G210), .B1(G237), .B2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G125), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(new_n224), .C1(new_n227), .C2(new_n230), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n241), .B2(new_n402), .ZN(new_n404));
  INV_X1    g218(.A(G224), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT7), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT8), .ZN(new_n411));
  INV_X1    g225(.A(G119), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G116), .ZN(new_n413));
  INV_X1    g227(.A(G116), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G119), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT89), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n248), .A2(new_n418), .A3(KEYINPUT5), .ZN(new_n419));
  INV_X1    g233(.A(G113), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n414), .A2(G119), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(new_n342), .A3(new_n255), .A4(new_n343), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n416), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n342), .A2(new_n343), .B1(new_n255), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n427), .B2(KEYINPUT90), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n255), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n371), .A2(new_n429), .A3(KEYINPUT90), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n411), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n408), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n403), .B(new_n432), .C1(new_n241), .C2(new_n402), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n409), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n409), .A2(new_n431), .A3(KEYINPUT91), .A4(new_n433), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n371), .A2(new_n429), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n350), .A2(new_n256), .A3(new_n352), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n410), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  INV_X1    g256(.A(new_n410), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT88), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n404), .A2(new_n406), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n403), .B(new_n407), .C1(new_n241), .C2(new_n402), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n442), .B(new_n443), .C1(KEYINPUT88), .C2(new_n445), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n324), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n401), .B1(new_n441), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(new_n324), .A3(new_n400), .A4(new_n452), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n399), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n261), .A2(G952), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(G234), .B2(G237), .ZN(new_n459));
  AOI211_X1 g273(.A(new_n324), .B(new_n261), .C1(G234), .C2(G237), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(G898), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n355), .A2(new_n356), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n260), .A2(new_n261), .A3(G214), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n260), .A2(new_n261), .A3(G214), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n467), .A2(new_n468), .B1(G143), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(KEYINPUT92), .A3(new_n466), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n195), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n218), .A2(new_n219), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n468), .B1(new_n473), .B2(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(G143), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G131), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G125), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n402), .A2(G140), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT16), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n402), .A2(KEYINPUT16), .A3(G140), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(G146), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n480), .A2(new_n481), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT19), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n222), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n478), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G113), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n331), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n476), .A2(KEYINPUT18), .A3(G131), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n485), .B(new_n222), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT18), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n470), .B(new_n471), .C1(new_n495), .C2(new_n195), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n493), .B(new_n494), .C1(new_n496), .C2(KEYINPUT93), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n476), .B1(KEYINPUT18), .B2(G131), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT94), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n493), .A2(new_n494), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n499), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(KEYINPUT93), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n492), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(G475), .A2(G902), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n472), .A2(new_n477), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n477), .A2(new_n510), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n482), .A2(new_n483), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n222), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n484), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n501), .A2(new_n506), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n508), .B(new_n509), .C1(new_n491), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT20), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n501), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n507), .B1(new_n522), .B2(new_n490), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n509), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n491), .A2(KEYINPUT95), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(KEYINPUT95), .A3(new_n491), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n324), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n519), .A2(new_n525), .B1(G475), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G122), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G116), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n329), .B1(new_n532), .B2(KEYINPUT14), .ZN(new_n533));
  XNOR2_X1  g347(.A(G116), .B(G122), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G143), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT97), .B1(new_n536), .B2(G128), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n225), .A3(G143), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n218), .A2(G128), .A3(new_n219), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n540), .A2(new_n541), .A3(new_n210), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n210), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n535), .B(KEYINPUT98), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n534), .B(G107), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n542), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n540), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n541), .A2(new_n551), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n541), .A2(KEYINPUT96), .A3(new_n551), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n550), .B1(new_n557), .B2(new_n189), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G217), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n395), .A2(new_n560), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n548), .A2(new_n558), .A3(new_n561), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n530), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n397), .A2(new_n464), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n560), .B1(G234), .B2(new_n324), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT79), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n412), .B2(G128), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT23), .B1(new_n225), .B2(G119), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n225), .A2(KEYINPUT79), .A3(G119), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT23), .A2(G119), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(G128), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n225), .A2(KEYINPUT78), .A3(KEYINPUT23), .A4(G119), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G110), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT81), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT81), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n580), .A2(new_n585), .A3(new_n589), .A4(new_n586), .ZN(new_n590));
  XOR2_X1   g404(.A(G119), .B(G128), .Z(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT24), .B(G110), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n485), .A2(new_n222), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n484), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n591), .A2(new_n592), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n580), .A2(new_n585), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(G110), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT80), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n600), .A2(new_n515), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n601), .B1(new_n600), .B2(new_n515), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT82), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT82), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n597), .B(new_n606), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n575), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n607), .A2(new_n575), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT25), .B1(new_n610), .B2(new_n324), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT25), .ZN(new_n612));
  NOR4_X1   g426(.A1(new_n608), .A2(new_n609), .A3(new_n612), .A4(G902), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n571), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n610), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n571), .A2(G902), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT83), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT84), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n322), .A2(new_n570), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  NAND2_X1  g438(.A1(new_n293), .A2(new_n324), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n625), .A2(G472), .B1(new_n294), .B2(new_n293), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n620), .B(KEYINPUT84), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n397), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n529), .A2(G475), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n517), .A2(new_n491), .ZN(new_n631));
  INV_X1    g445(.A(new_n509), .ZN(new_n632));
  NOR4_X1   g446(.A1(new_n631), .A2(KEYINPUT20), .A3(new_n507), .A4(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n524), .B1(new_n523), .B2(new_n509), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n566), .A2(G902), .ZN(new_n636));
  INV_X1    g450(.A(new_n564), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n561), .B1(new_n548), .B2(new_n558), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n637), .A2(KEYINPUT33), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n563), .B2(new_n564), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(G478), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n565), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n324), .B1(new_n637), .B2(new_n638), .ZN(new_n646));
  INV_X1    g460(.A(new_n644), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT100), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n642), .B(KEYINPUT101), .C1(new_n645), .C2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n643), .B1(new_n565), .B2(new_n644), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT101), .B1(new_n653), .B2(new_n642), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n635), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT102), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n635), .B(new_n657), .C1(new_n650), .C2(new_n654), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n464), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n629), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT34), .B(G104), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(new_n568), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n530), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n464), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n629), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n625), .A2(G472), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n604), .B(KEYINPUT103), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n575), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n617), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n614), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n669), .A2(new_n295), .A3(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n570), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT105), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n679), .B(new_n681), .ZN(G12));
  NAND4_X1  g496(.A1(new_n394), .A2(new_n675), .A3(new_n457), .A4(new_n396), .ZN(new_n683));
  INV_X1    g497(.A(new_n459), .ZN(new_n684));
  INV_X1    g498(.A(new_n460), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n684), .B1(new_n685), .B2(G900), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n530), .A2(new_n663), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n322), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  AND2_X1   g504(.A1(new_n454), .A2(new_n456), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n399), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n686), .B(KEYINPUT39), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n394), .A2(new_n396), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n530), .A2(new_n568), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n693), .A2(new_n696), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n308), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n265), .B1(new_n700), .B2(new_n258), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n303), .B2(new_n269), .ZN(new_n702));
  OAI21_X1  g516(.A(G472), .B1(new_n702), .B2(G902), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n297), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n321), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT77), .B1(new_n293), .B2(new_n298), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n699), .A2(new_n709), .A3(new_n675), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n465), .ZN(G45));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n635), .B(new_n686), .C1(new_n650), .C2(new_n654), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n683), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n712), .B1(new_n322), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n322), .A2(new_n714), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  AOI22_X1  g533(.A1(new_n296), .A2(new_n295), .B1(new_n319), .B2(G472), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n628), .B1(new_n707), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n382), .A2(new_n386), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n396), .A3(new_n387), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n659), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT107), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n726), .B(new_n728), .ZN(G15));
  NAND4_X1  g543(.A1(new_n322), .A2(new_n725), .A3(new_n622), .A4(new_n665), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT108), .B(G116), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G18));
  NAND4_X1  g546(.A1(new_n723), .A2(new_n463), .A3(new_n396), .A4(new_n387), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n675), .A2(new_n457), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n733), .A2(new_n734), .A3(new_n569), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n322), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n669), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n625), .A2(KEYINPUT110), .A3(G472), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n698), .A2(new_n457), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n733), .ZN(new_n743));
  INV_X1    g557(.A(new_n620), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n309), .A2(new_n265), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n282), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n282), .A2(new_n745), .A3(KEYINPUT109), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n292), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n294), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n741), .A2(new_n743), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NOR3_X1   g567(.A1(new_n713), .A2(new_n734), .A3(new_n724), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n741), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  AND3_X1   g570(.A1(new_n454), .A2(new_n398), .A3(new_n456), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n394), .A2(new_n757), .A3(new_n396), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n394), .A2(new_n757), .A3(new_n760), .A4(new_n396), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n713), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n721), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n759), .A2(new_n763), .A3(new_n761), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n297), .A2(new_n320), .A3(new_n305), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(new_n744), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n768), .B2(new_n744), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT42), .B(new_n767), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  INV_X1    g588(.A(new_n687), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n721), .A2(new_n762), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n779));
  INV_X1    g593(.A(new_n391), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n327), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n781), .B2(new_n389), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n782), .B2(new_n323), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n780), .A2(new_n327), .B1(new_n383), .B2(new_n388), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT45), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT113), .B(G469), .C1(new_n784), .C2(KEYINPUT45), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n393), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n393), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n387), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n396), .ZN(new_n793));
  INV_X1    g607(.A(new_n694), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n778), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(KEYINPUT114), .A3(new_n396), .A4(new_n694), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n530), .B1(new_n650), .B2(new_n654), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT43), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT43), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n627), .A2(new_n675), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n802), .B2(new_n803), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n757), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n795), .A2(new_n796), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  INV_X1    g623(.A(new_n757), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n322), .A2(new_n622), .A3(new_n713), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n396), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT47), .B1(new_n792), .B2(new_n396), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  AOI22_X1  g630(.A1(new_n739), .A2(new_n740), .B1(new_n294), .B2(new_n750), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n675), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n724), .A2(new_n810), .A3(new_n684), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n800), .A2(new_n801), .A3(new_n819), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n818), .A2(new_n820), .A3(KEYINPUT121), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT121), .B1(new_n818), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n709), .A2(new_n622), .A3(new_n819), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n635), .A2(new_n650), .A3(new_n654), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n800), .A2(new_n459), .A3(new_n801), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n744), .A3(new_n725), .A4(new_n817), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n692), .A2(new_n399), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n817), .A2(new_n744), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n800), .A2(new_n459), .A3(new_n801), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n833), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n725), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n829), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n723), .A2(new_n387), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n396), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n813), .A2(new_n814), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n757), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n828), .B(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n656), .A2(new_n658), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n458), .B1(new_n824), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n457), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n832), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n768), .A2(new_n744), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT112), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n768), .A2(new_n769), .A3(new_n744), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(new_n820), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT47), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n793), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n812), .C1(new_n396), .C2(new_n841), .ZN(new_n861));
  INV_X1    g675(.A(new_n844), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n827), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n834), .A2(KEYINPUT120), .A3(new_n839), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT120), .B1(new_n834), .B2(new_n839), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n845), .B(new_n858), .C1(new_n867), .C2(KEYINPUT51), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n726), .A2(new_n730), .A3(new_n736), .A4(new_n752), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n773), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n322), .A2(new_n712), .A3(new_n714), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n689), .B(new_n755), .C1(new_n872), .C2(new_n715), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n686), .B(KEYINPUT117), .Z(new_n874));
  NOR3_X1   g688(.A1(new_n742), .A2(new_n397), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n675), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n708), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n871), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n817), .A2(new_n754), .B1(new_n322), .B2(new_n688), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n718), .A2(KEYINPUT52), .A3(new_n880), .A4(new_n877), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n870), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n397), .A2(new_n464), .ZN(new_n883));
  INV_X1    g697(.A(new_n655), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n622), .A2(new_n883), .A3(new_n626), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n623), .A2(new_n885), .A3(KEYINPUT116), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n679), .A2(new_n886), .A3(new_n666), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n767), .A2(new_n817), .A3(new_n675), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n675), .A2(new_n686), .ZN(new_n889));
  INV_X1    g703(.A(new_n569), .ZN(new_n890));
  INV_X1    g704(.A(new_n758), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n322), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n776), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT116), .B1(new_n623), .B2(new_n885), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n887), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n879), .A2(new_n881), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n767), .A2(KEYINPUT42), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n898), .A2(new_n853), .B1(new_n764), .B2(new_n765), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n726), .A2(new_n730), .A3(new_n752), .A4(new_n736), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n879), .B2(new_n881), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n869), .A2(new_n773), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT119), .B1(new_n899), .B2(new_n900), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n895), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n905), .A2(new_n914), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n868), .A2(new_n915), .B1(G952), .B2(G953), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n692), .A2(new_n744), .A3(new_n398), .A4(new_n396), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n841), .B(KEYINPUT49), .ZN(new_n918));
  OR4_X1    g732(.A1(new_n708), .A2(new_n917), .A3(new_n918), .A4(new_n797), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(G75));
  NAND2_X1  g734(.A1(new_n906), .A2(new_n913), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(G210), .A3(G902), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n447), .A2(new_n451), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n450), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n261), .A2(G952), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G51));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  INV_X1    g745(.A(new_n787), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n931), .A2(new_n921), .A3(G902), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n324), .B1(new_n906), .B2(new_n913), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n393), .B(KEYINPUT57), .Z(new_n937));
  AND3_X1   g751(.A1(new_n906), .A2(new_n907), .A3(new_n913), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n907), .B1(new_n906), .B2(new_n913), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n722), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n929), .B1(new_n936), .B2(new_n942), .ZN(G54));
  NAND3_X1  g757(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n631), .B2(new_n507), .ZN(new_n945));
  INV_X1    g759(.A(new_n929), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .A4(new_n523), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G60));
  NOR2_X1   g762(.A1(new_n639), .A2(new_n641), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT59), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n950), .B(new_n952), .C1(new_n938), .C2(new_n939), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n946), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n915), .B2(new_n952), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G63));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n906), .B2(new_n913), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n672), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n946), .B1(new_n960), .B2(new_n610), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n960), .A2(new_n610), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n461), .B2(new_n405), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n623), .A2(new_n885), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT116), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n666), .A3(new_n679), .A4(new_n886), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n261), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n974), .B2(new_n261), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n968), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  INV_X1    g796(.A(G898), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n924), .B1(new_n983), .B2(G953), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n980), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n980), .B2(new_n982), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n270), .A2(new_n279), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(new_n486), .Z(new_n990));
  NOR2_X1   g804(.A1(new_n854), .A2(new_n742), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n795), .A2(new_n796), .A3(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n776), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n899), .A2(new_n993), .A3(new_n873), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n808), .A2(new_n992), .A3(new_n815), .A4(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n988), .B(new_n990), .C1(new_n995), .C2(G953), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n808), .A2(new_n815), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n710), .A2(new_n873), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n710), .B2(new_n873), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n810), .B(new_n695), .C1(new_n655), .C2(new_n664), .ZN(new_n1001));
  AOI22_X1  g815(.A1(new_n999), .A2(new_n1000), .B1(new_n721), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(G953), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n990), .B(KEYINPUT125), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n995), .B2(new_n974), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n315), .A2(new_n265), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT127), .Z(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n316), .A2(new_n281), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1009), .B(new_n1014), .C1(new_n896), .C2(new_n904), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1013), .A2(new_n946), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n997), .A2(new_n973), .A3(new_n1002), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT126), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1017), .A2(new_n1018), .A3(new_n1009), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n315), .A2(new_n265), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1017), .A2(new_n1009), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(KEYINPUT126), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1016), .B1(new_n1019), .B2(new_n1022), .ZN(G57));
endmodule


