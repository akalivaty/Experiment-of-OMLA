//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n204));
  INV_X1    g0004(.A(G87), .ZN(new_n205));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT64), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n211), .B(new_n212), .C1(G77), .C2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n203), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n223), .A2(new_n226), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n217), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NOR2_X1   g0048(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT13), .ZN(new_n250));
  AND2_X1   g0050(.A1(G232), .A2(G1698), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  OAI211_X1 g0058(.A(G226), .B(new_n258), .C1(new_n252), .C2(new_n253), .ZN(new_n259));
  OAI211_X1 g0059(.A(KEYINPUT72), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n256), .A2(new_n257), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n215), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT73), .ZN(new_n273));
  AND4_X1   g0073(.A1(new_n250), .A2(new_n265), .A3(new_n270), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n269), .B1(new_n261), .B2(new_n264), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n250), .B1(new_n275), .B2(new_n273), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n249), .B1(new_n277), .B2(G179), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n265), .A2(new_n270), .A3(new_n273), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n275), .A2(new_n250), .A3(new_n273), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n280), .B1(new_n284), .B2(G169), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  AOI211_X1 g0086(.A(new_n286), .B(new_n279), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n278), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT76), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT67), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n293), .A2(new_n266), .A3(G13), .A4(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n214), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(KEYINPUT12), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT12), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(KEYINPUT74), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(KEYINPUT74), .B2(new_n299), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n229), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n292), .B2(new_n294), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n266), .A2(KEYINPUT68), .A3(G20), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT68), .B1(new_n266), .B2(G20), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(G68), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n228), .A2(G33), .A3(G77), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G20), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n309), .B1(new_n228), .B2(G68), .C1(new_n311), .C2(new_n219), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n303), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT11), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n301), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n278), .B(KEYINPUT76), .C1(new_n285), .C2(new_n287), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n290), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n284), .A2(G200), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n277), .A2(G190), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT77), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT3), .B(G33), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(G20), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n252), .A2(new_n253), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n214), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G58), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n214), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G58), .A2(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n310), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n324), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT7), .B1(new_n326), .B2(G20), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n328), .A2(new_n325), .A3(new_n228), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(G68), .ZN(new_n340));
  INV_X1    g0140(.A(new_n336), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n342), .A3(new_n303), .ZN(new_n343));
  INV_X1    g0143(.A(new_n303), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n295), .A2(new_n307), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT8), .A2(G58), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT8), .A2(G58), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT79), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n292), .B2(new_n294), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n346), .A2(new_n347), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n304), .B2(new_n307), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT79), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT80), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n353), .B2(new_n356), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n343), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G223), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n258), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n326), .B(new_n362), .C1(G226), .C2(new_n258), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n263), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n272), .ZN(new_n366));
  INV_X1    g0166(.A(G232), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n268), .A2(new_n367), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G179), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n286), .B2(new_n369), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT18), .B1(new_n360), .B2(new_n371), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n343), .B(new_n377), .C1(new_n358), .C2(new_n359), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n369), .A2(G190), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n343), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n350), .B1(new_n349), .B2(new_n352), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n355), .A2(KEYINPUT79), .A3(new_n351), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT80), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(KEYINPUT81), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n387), .A2(new_n390), .A3(new_n379), .A4(new_n377), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT15), .B(G87), .Z(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(new_n228), .A3(G33), .ZN(new_n394));
  INV_X1    g0194(.A(G77), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n310), .B(KEYINPUT69), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n394), .B1(new_n228), .B2(new_n395), .C1(new_n354), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n303), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n296), .A2(new_n395), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n395), .C2(new_n345), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G238), .A2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n326), .B(new_n401), .C1(new_n367), .C2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n264), .C1(G107), .C2(new_n326), .ZN(new_n403));
  INV_X1    g0203(.A(new_n268), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G244), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n272), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n400), .B1(G190), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n376), .B2(new_n407), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n374), .A2(new_n392), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n323), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G33), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n354), .A2(G20), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G150), .ZN(new_n414));
  NOR3_X1   g0214(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n414), .A2(new_n311), .B1(new_n415), .B2(new_n228), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n303), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n296), .A2(new_n219), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n219), .C2(new_n345), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT70), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT9), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n424), .A2(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n258), .A2(G222), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n326), .B(new_n426), .C1(new_n361), .C2(new_n258), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n264), .C1(G77), .C2(new_n326), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n272), .C1(new_n220), .C2(new_n268), .ZN(new_n429));
  INV_X1    g0229(.A(G190), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n425), .B(new_n431), .C1(G200), .C2(new_n429), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n424), .A2(KEYINPUT10), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n423), .B(new_n432), .C1(new_n424), .C2(KEYINPUT10), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(new_n286), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n419), .C1(G179), .C2(new_n429), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n406), .A2(new_n286), .ZN(new_n440));
  INV_X1    g0240(.A(G179), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n407), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n400), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n411), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n228), .C1(G33), .C2(new_n207), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n302), .A2(new_n229), .B1(G20), .B2(new_n216), .ZN(new_n450));
  AOI21_X1  g0250(.A(G20), .B1(new_n412), .B2(G97), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT87), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n447), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n449), .A2(new_n453), .A3(KEYINPUT20), .A4(new_n450), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n296), .A2(new_n216), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n266), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n304), .A2(G116), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G264), .A2(G1698), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n326), .B(new_n463), .C1(new_n208), .C2(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n264), .C1(G303), .C2(new_n326), .ZN(new_n465));
  INV_X1    g0265(.A(G41), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n266), .B(G45), .C1(new_n466), .C2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  OAI211_X1 g0269(.A(G270), .B(new_n263), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(KEYINPUT82), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(G274), .B1(new_n468), .B2(G41), .ZN(new_n478));
  INV_X1    g0278(.A(new_n229), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n262), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n477), .A2(KEYINPUT83), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT83), .B1(new_n477), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n465), .B(new_n470), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n462), .A2(G169), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT88), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n462), .A2(new_n483), .A3(new_n487), .A4(G169), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT89), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n483), .A2(KEYINPUT21), .A3(G169), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n483), .A2(new_n441), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n462), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n485), .A2(KEYINPUT89), .A3(new_n486), .A4(new_n488), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n483), .A2(G200), .ZN(new_n496));
  INV_X1    g0296(.A(new_n462), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n497), .C1(new_n430), .C2(new_n483), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n491), .A2(new_n494), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G20), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT23), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n228), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n326), .A2(new_n506), .A3(new_n228), .A4(G87), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n303), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n304), .A2(new_n460), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n501), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n296), .A2(new_n501), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT25), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n507), .ZN(new_n523));
  INV_X1    g0323(.A(new_n503), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n510), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT24), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n515), .B1(new_n528), .B2(new_n303), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(KEYINPUT90), .A3(new_n519), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n467), .A2(KEYINPUT82), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n480), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n477), .A2(KEYINPUT83), .A3(new_n480), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n206), .A2(new_n258), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n208), .A2(G1698), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n252), .C2(new_n253), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n263), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G264), .B(new_n263), .C1(new_n467), .C2(new_n469), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n537), .A2(G179), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n481), .B2(new_n482), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(KEYINPUT91), .A3(G169), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT91), .B1(new_n547), .B2(G169), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n522), .A2(new_n530), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT92), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n547), .A2(new_n553), .A3(new_n376), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n547), .B2(new_n376), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n545), .B(new_n430), .C1(new_n481), .C2(new_n482), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n520), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n295), .A2(G97), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n514), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n501), .B1(new_n327), .B2(new_n329), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n311), .A2(new_n395), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT6), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n207), .A2(new_n501), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n501), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n228), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n561), .B(new_n563), .C1(new_n572), .C2(new_n344), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(new_n263), .C1(new_n467), .C2(new_n469), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n326), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n576));
  OAI21_X1  g0376(.A(G244), .B1(new_n252), .B2(new_n253), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n579), .A3(new_n447), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n326), .A2(G250), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n258), .B1(new_n581), .B2(KEYINPUT4), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n264), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n537), .A2(new_n575), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n574), .B(new_n585), .C1(new_n430), .C2(new_n584), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n286), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n537), .A2(new_n583), .A3(new_n441), .A4(new_n575), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n573), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n552), .A2(new_n559), .A3(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G238), .B(new_n258), .C1(new_n252), .C2(new_n253), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT84), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n326), .A2(KEYINPUT84), .A3(G238), .A4(new_n258), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n326), .A2(G244), .A3(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n264), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n473), .A2(new_n271), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n206), .B1(new_n472), .B2(G1), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n263), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT85), .ZN(new_n604));
  INV_X1    g0404(.A(new_n602), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n598), .B2(new_n264), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n286), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n599), .B2(new_n602), .ZN(new_n610));
  AOI211_X1 g0410(.A(KEYINPUT85), .B(new_n605), .C1(new_n598), .C2(new_n264), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n441), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n326), .A2(new_n228), .A3(G68), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n568), .A2(new_n205), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n257), .A2(new_n228), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(KEYINPUT19), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n257), .B2(G20), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n303), .ZN(new_n620));
  INV_X1    g0420(.A(new_n393), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n296), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT86), .B1(new_n620), .B2(new_n622), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n624), .A2(new_n625), .B1(new_n514), .B2(new_n621), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n609), .A2(new_n612), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n604), .A2(G200), .A3(new_n608), .ZN(new_n628));
  OAI21_X1  g0428(.A(G190), .B1(new_n610), .B2(new_n611), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(new_n622), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n623), .B1(G87), .B2(new_n562), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n500), .A2(new_n591), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n446), .A2(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n321), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n317), .B1(new_n443), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n392), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n372), .A2(new_n373), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n435), .B(new_n436), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n438), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT93), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n603), .A2(new_n645), .A3(new_n286), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT93), .B1(new_n606), .B2(G169), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n612), .A3(new_n626), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n603), .A2(G200), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n629), .A2(new_n633), .A3(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n649), .B(new_n651), .C1(new_n558), .C2(new_n520), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n590), .ZN(new_n653));
  INV_X1    g0453(.A(new_n550), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n546), .A3(new_n548), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n520), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n491), .A2(new_n494), .A3(new_n656), .A4(new_n495), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n587), .A2(new_n573), .A3(new_n588), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n627), .A2(new_n634), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n649), .A2(new_n659), .A3(new_n651), .A4(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n649), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n644), .B1(new_n446), .B2(new_n665), .ZN(G369));
  NAND3_X1  g0466(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n266), .A2(new_n228), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n462), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n499), .B(KEYINPUT94), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT90), .B1(new_n529), .B2(new_n519), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n344), .B1(new_n526), .B2(new_n527), .ZN(new_n680));
  NOR4_X1   g0480(.A1(new_n680), .A2(new_n521), .A3(new_n518), .A4(new_n515), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n673), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT95), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n655), .B1(new_n679), .B2(new_n681), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n683), .B(new_n684), .C1(new_n520), .C2(new_n558), .ZN(new_n685));
  INV_X1    g0485(.A(new_n673), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n656), .A2(new_n673), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n667), .A2(new_n686), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n224), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n568), .A2(new_n205), .A3(new_n216), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(new_n266), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n699));
  INV_X1    g0499(.A(new_n695), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n698), .B(new_n699), .C1(new_n227), .C2(new_n700), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT97), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n665), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n684), .A2(new_n494), .A3(new_n491), .A4(new_n495), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n653), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT99), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n649), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n649), .A2(new_n659), .A3(new_n651), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(KEYINPUT26), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(KEYINPUT99), .A3(new_n653), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n686), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n704), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n500), .A2(new_n591), .A3(new_n636), .A4(new_n686), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n604), .A2(new_n608), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n537), .A2(new_n583), .A3(new_n545), .A4(new_n575), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n493), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n493), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n584), .A2(new_n547), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT98), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT98), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n584), .A2(new_n726), .A3(new_n547), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n441), .A3(new_n483), .A4(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n722), .B(new_n723), .C1(new_n728), .C2(new_n606), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n673), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n716), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n715), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT100), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n703), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(G13), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n266), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n695), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n678), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n677), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n677), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n228), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n441), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n376), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G329), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n757), .A2(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n441), .A2(new_n376), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n751), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n755), .B(new_n762), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n228), .A2(new_n430), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n752), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G322), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n763), .A2(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G326), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n228), .B1(new_n759), .B2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G294), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n767), .A2(new_n771), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n768), .A2(new_n756), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n328), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT102), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n764), .A2(new_n214), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n772), .A2(new_n219), .B1(new_n753), .B2(new_n395), .ZN(new_n784));
  INV_X1    g0584(.A(new_n757), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G107), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n760), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(KEYINPUT32), .A3(G159), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT32), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n760), .B2(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n788), .A2(new_n791), .B1(G58), .B2(new_n770), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n776), .A2(G97), .ZN(new_n793));
  INV_X1    g0593(.A(new_n779), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n328), .B1(new_n794), .B2(G87), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n786), .A2(new_n792), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n778), .A2(new_n782), .B1(new_n783), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n229), .B1(G20), .B2(new_n286), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n748), .A2(new_n798), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n694), .A2(new_n326), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(G45), .B2(new_n227), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT101), .Z(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n244), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n694), .A2(new_n328), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G355), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G116), .B2(new_n224), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n800), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n750), .A2(new_n799), .A3(new_n808), .A4(new_n743), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n745), .A2(new_n809), .ZN(G396));
  XNOR2_X1  g0610(.A(new_n443), .B(KEYINPUT105), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n409), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n686), .B(new_n813), .C1(new_n658), .C2(new_n664), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n400), .A2(new_n673), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n443), .B2(new_n686), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n663), .A2(new_n649), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n653), .A2(new_n657), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n673), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n814), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(new_n735), .ZN(new_n824));
  INV_X1    g0624(.A(new_n743), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n735), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n793), .B1(new_n501), .B2(new_n779), .C1(new_n754), .C2(new_n760), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n328), .B1(new_n769), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n205), .A2(new_n757), .B1(new_n753), .B2(new_n216), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n758), .B2(new_n764), .C1(new_n780), .C2(new_n772), .ZN(new_n833));
  INV_X1    g0633(.A(new_n753), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G143), .A2(new_n770), .B1(new_n834), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n836), .B2(new_n772), .C1(new_n414), .C2(new_n764), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT104), .ZN(new_n838));
  XOR2_X1   g0638(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n839));
  XNOR2_X1  g0639(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n840), .B1(new_n331), .B2(new_n775), .C1(new_n214), .C2(new_n757), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n326), .B1(new_n760), .B2(new_n842), .C1(new_n219), .C2(new_n779), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n833), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n798), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n813), .A2(new_n815), .B1(new_n444), .B2(new_n673), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n746), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n798), .A2(new_n746), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n395), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n845), .A2(new_n743), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n827), .A2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT109), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n392), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n381), .A2(new_n391), .A3(KEYINPUT109), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n374), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n387), .A2(new_n671), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n671), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n360), .B1(new_n371), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n385), .A2(new_n386), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n860), .A2(new_n343), .A3(new_n379), .A4(new_n377), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n342), .A2(new_n303), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT16), .B1(new_n340), .B2(new_n341), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n383), .A2(new_n384), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n371), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n378), .B2(new_n380), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT108), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n858), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT107), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT107), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n868), .A2(new_n874), .A3(new_n858), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT108), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n861), .A2(new_n878), .A3(new_n869), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n871), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n865), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n877), .B1(new_n374), .B2(new_n392), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT40), .B1(new_n864), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n316), .ZN(new_n886));
  OAI21_X1  g0686(.A(G169), .B1(new_n274), .B2(new_n276), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n279), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n284), .A2(G169), .A3(new_n280), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT76), .B1(new_n890), .B2(new_n278), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n315), .B(new_n673), .C1(new_n892), .C2(new_n639), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n315), .A2(new_n673), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n317), .A2(new_n321), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n846), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n734), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n885), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n895), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT110), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n734), .A3(new_n901), .A4(new_n817), .ZN(new_n902));
  INV_X1    g0702(.A(new_n865), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n861), .A2(new_n878), .A3(new_n869), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n878), .B1(new_n861), .B2(new_n869), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n904), .A2(new_n905), .A3(new_n876), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n374), .A2(new_n392), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n876), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n901), .B1(new_n896), .B2(new_n734), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n899), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT111), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT111), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n899), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n898), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n411), .A2(new_n445), .A3(new_n734), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT112), .Z(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G330), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n644), .B1(new_n446), .B2(new_n715), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n864), .B2(new_n884), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n892), .A2(new_n315), .A3(new_n686), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT39), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n811), .A2(new_n673), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n814), .A2(new_n933), .B1(new_n895), .B2(new_n893), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n913), .B1(new_n642), .B2(new_n671), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n925), .B(new_n936), .Z(new_n937));
  XNOR2_X1  g0737(.A(new_n924), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n266), .B2(new_n740), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n569), .A2(new_n570), .ZN(new_n940));
  OAI211_X1 g0740(.A(G20), .B(new_n479), .C1(new_n940), .C2(KEYINPUT35), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n216), .B(new_n941), .C1(KEYINPUT35), .C2(new_n940), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT36), .Z(new_n943));
  NOR3_X1   g0743(.A1(new_n332), .A2(new_n227), .A3(new_n395), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT106), .Z(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(G50), .B2(new_n214), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n739), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n939), .A2(new_n943), .A3(new_n947), .ZN(G367));
  OAI211_X1 g0748(.A(new_n586), .B(new_n589), .C1(new_n574), .C2(new_n686), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n589), .B1(new_n949), .B2(new_n684), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n686), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT42), .B1(new_n692), .B2(new_n949), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n649), .A2(new_n633), .A3(new_n686), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n649), .B(new_n651), .C1(new_n633), .C2(new_n686), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n659), .A2(new_n673), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n688), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n959), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n695), .B(KEYINPUT41), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n692), .A2(new_n690), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n962), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n692), .A2(new_n690), .A3(new_n961), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT45), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n688), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT115), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT115), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n972), .A2(new_n974), .A3(new_n978), .A4(new_n688), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n678), .A2(new_n687), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n688), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(new_n691), .Z(new_n983));
  XOR2_X1   g0783(.A(new_n688), .B(KEYINPUT114), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n975), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n983), .A3(new_n737), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n968), .B1(new_n986), .B2(new_n737), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n966), .B1(new_n987), .B2(new_n742), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n328), .B1(new_n775), .B2(new_n501), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n757), .A2(new_n207), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G317), .B2(new_n787), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n758), .B2(new_n753), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n989), .B(new_n992), .C1(G303), .C2(new_n770), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT116), .B(G311), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n773), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n794), .A2(G116), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n765), .A2(G294), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n993), .A2(new_n995), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n326), .B1(new_n769), .B2(new_n414), .C1(new_n331), .C2(new_n779), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n773), .A2(G143), .B1(new_n776), .B2(G68), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n836), .B2(new_n760), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G159), .B2(new_n765), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n785), .A2(G77), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n219), .C2(new_n753), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n999), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n798), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n955), .A2(new_n748), .A3(new_n956), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n801), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n800), .B1(new_n224), .B2(new_n621), .C1(new_n239), .C2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n743), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n988), .A2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n983), .A2(new_n737), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n983), .A2(new_n737), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n695), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n621), .A2(new_n775), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G50), .B2(new_n770), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n395), .B2(new_n779), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n326), .B1(new_n772), .B2(new_n790), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n990), .B1(G68), .B2(new_n834), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n354), .B2(new_n764), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n414), .B2(new_n760), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G322), .A2(new_n773), .B1(new_n770), .B2(G317), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n765), .A2(new_n994), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n780), .C2(new_n753), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n758), .B2(new_n775), .C1(new_n829), .C2(new_n779), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n785), .A2(G116), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n787), .A2(G326), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1031), .A2(new_n328), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1024), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n236), .A2(new_n472), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n801), .B1(new_n696), .B2(new_n805), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n348), .A2(new_n219), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n214), .A2(new_n395), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1040), .A2(G45), .A3(new_n1041), .A4(new_n696), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1038), .A2(new_n1042), .B1(G107), .B2(new_n224), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1036), .A2(new_n798), .B1(new_n800), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n743), .B(new_n1044), .C1(new_n687), .C2(new_n749), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT117), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n983), .C2(new_n742), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1016), .A2(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n975), .A2(new_n976), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n980), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(new_n741), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n800), .B1(new_n207), .B2(new_n224), .C1(new_n247), .C2(new_n1010), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n961), .B2(new_n749), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G317), .A2(new_n773), .B1(new_n770), .B2(G311), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G116), .B2(new_n776), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n834), .A2(G294), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G107), .A2(new_n785), .B1(new_n787), .B2(G322), .ZN(new_n1060));
  AND4_X1   g0860(.A1(new_n328), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n758), .B2(new_n779), .C1(new_n780), .C2(new_n764), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n772), .A2(new_n414), .B1(new_n769), .B2(new_n790), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n348), .B2(new_n834), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n219), .B2(new_n764), .C1(new_n395), .C2(new_n775), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n328), .B1(new_n787), .B2(G143), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n214), .B2(new_n779), .C1(new_n205), .C2(new_n757), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT118), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1062), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n825), .B(new_n1055), .C1(new_n798), .C2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1053), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1052), .A2(new_n1015), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n695), .A3(new_n986), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(KEYINPUT119), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n734), .A2(G330), .A3(new_n817), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n317), .A2(new_n321), .A3(new_n894), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n894), .B1(new_n317), .B2(new_n321), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1076), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(G330), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n732), .A2(new_n733), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1082), .B1(new_n1083), .B2(new_n716), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1084), .A2(KEYINPUT119), .A3(new_n817), .A4(new_n900), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n735), .A2(KEYINPUT120), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT120), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n734), .A2(new_n1088), .A3(G330), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n817), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1080), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n713), .A2(new_n686), .A3(new_n813), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n933), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1086), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1084), .A2(new_n817), .A3(new_n900), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n932), .B1(new_n822), .B2(new_n813), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n411), .A2(G330), .A3(new_n445), .A4(new_n734), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n644), .C1(new_n446), .C2(new_n715), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n928), .B1(new_n1099), .B2(new_n1080), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n381), .A2(new_n391), .A3(KEYINPUT109), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT109), .B1(new_n381), .B2(new_n391), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n642), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n856), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n863), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n883), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT39), .B1(new_n1113), .B2(new_n911), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1080), .B1(new_n1092), .B2(new_n933), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n928), .B1(new_n864), .B2(new_n884), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1116), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1093), .B2(new_n900), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n673), .B(new_n812), .C1(new_n820), .C2(new_n821), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n900), .B1(new_n1122), .B2(new_n932), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n927), .A2(new_n930), .B1(new_n1123), .B2(new_n928), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1096), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1106), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1126), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1093), .B1(new_n1090), .B2(new_n1080), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1129), .A2(new_n1086), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1104), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1132), .A3(new_n695), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n742), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n746), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n848), .A2(new_n354), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n753), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n779), .A2(new_n414), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n776), .A2(G159), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n326), .B1(new_n769), .B2(new_n842), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G125), .B2(new_n787), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n773), .A2(G128), .B1(new_n785), .B2(G50), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1138), .B(new_n1145), .C1(G137), .C2(new_n765), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n328), .B1(new_n764), .B2(new_n501), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n779), .A2(new_n205), .B1(new_n757), .B2(new_n214), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(G77), .C2(new_n776), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G97), .A2(new_n834), .B1(new_n787), .B2(G294), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n758), .C2(new_n772), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G116), .B2(new_n770), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n798), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1135), .A2(new_n743), .A3(new_n1136), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1133), .A2(new_n1134), .A3(new_n1154), .ZN(G378));
  OAI21_X1  g0955(.A(new_n1105), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n439), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n435), .A2(new_n436), .A3(new_n438), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n421), .B2(new_n671), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n421), .A2(new_n671), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n931), .A2(new_n1165), .A3(new_n935), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n931), .B2(new_n935), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n920), .A2(G330), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n898), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n919), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n817), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n716), .A2(new_n732), .A3(new_n733), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT110), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n913), .A3(new_n902), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n918), .B1(new_n1175), .B2(new_n899), .ZN(new_n1176));
  OAI211_X1 g0976(.A(G330), .B(new_n1170), .C1(new_n1171), .C2(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1156), .A2(KEYINPUT57), .A3(new_n1169), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n695), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT121), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1168), .B1(new_n920), .B2(G330), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(new_n1169), .A3(KEYINPUT121), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1156), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1181), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1165), .A2(new_n746), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n395), .A2(new_n779), .B1(new_n769), .B2(new_n501), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G41), .B(new_n1192), .C1(G68), .C2(new_n776), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n326), .B1(new_n785), .B2(G58), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n834), .A2(new_n393), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n765), .A2(G97), .B1(new_n787), .B2(G283), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G116), .B2(new_n773), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT58), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n219), .B1(new_n252), .B2(G41), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n773), .A2(G125), .ZN(new_n1201));
  INV_X1    g1001(.A(G128), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n769), .A2(new_n1202), .B1(new_n753), .B2(new_n836), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n779), .A2(new_n1137), .B1(new_n775), .B2(new_n414), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n764), .A2(new_n842), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G33), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G41), .B1(new_n787), .B2(G124), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n790), .C2(new_n757), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1200), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n798), .B1(new_n1199), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n848), .A2(new_n219), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1191), .A2(new_n743), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1179), .A2(new_n1169), .A3(KEYINPUT121), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT121), .B1(new_n1179), .B2(new_n1169), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1219), .B2(new_n742), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1190), .A2(new_n1220), .ZN(G375));
  INV_X1    g1021(.A(new_n798), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n772), .A2(new_n842), .B1(new_n764), .B2(new_n1137), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G137), .B2(new_n770), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT123), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n326), .B1(new_n757), .B2(new_n331), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1202), .A2(new_n760), .B1(new_n775), .B2(new_n219), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n414), .B2(new_n753), .C1(new_n790), .C2(new_n779), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1004), .B1(new_n829), .B2(new_n772), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n328), .B1(new_n753), .B2(new_n501), .C1(new_n207), .C2(new_n779), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n760), .A2(new_n780), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1017), .A4(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n216), .B2(new_n764), .C1(new_n758), .C2(new_n769), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1222), .B1(new_n1229), .B2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n825), .B(new_n1235), .C1(new_n214), .C2(new_n848), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n900), .A2(new_n747), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT122), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1102), .A2(new_n742), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1095), .A2(new_n1104), .A3(new_n1101), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n967), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1239), .B1(new_n1241), .B2(new_n1131), .ZN(G381));
  NAND4_X1  g1042(.A1(new_n988), .A2(new_n1012), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1243));
  INV_X1    g1043(.A(G396), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1016), .A2(new_n1244), .A3(new_n1049), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1243), .A2(G384), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G375), .A2(G378), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(G407));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1246), .B2(new_n672), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(G213), .ZN(G409));
  NAND2_X1  g1050(.A1(G387), .A2(G390), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1245), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1244), .B1(new_n1016), .B2(new_n1049), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT127), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1253), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT127), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1245), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1251), .A2(new_n1258), .A3(new_n1243), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1251), .A2(new_n1243), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1257), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G343), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1156), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1220), .C1(new_n1265), .C2(new_n1181), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1186), .A2(new_n967), .A3(new_n1156), .A4(new_n1187), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1179), .A2(new_n1169), .A3(new_n742), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1215), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G378), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1264), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n827), .A2(KEYINPUT126), .A3(new_n850), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1240), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n695), .A3(new_n1106), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1240), .B2(new_n1274), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1239), .B(new_n1273), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G384), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1240), .A2(new_n1274), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT60), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1285), .A2(new_n695), .A3(new_n1106), .A4(new_n1276), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1239), .A3(new_n1281), .A4(new_n1273), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1186), .A2(new_n742), .A3(new_n1187), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1215), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1189), .A2(new_n1270), .A3(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT124), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1264), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1266), .A2(new_n1299), .A3(new_n1271), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1264), .A2(G2897), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1288), .B(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1290), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1297), .A2(new_n1298), .A3(new_n1288), .A4(new_n1300), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1262), .B(new_n1292), .C1(new_n1304), .C2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1261), .B1(new_n1251), .B2(new_n1243), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1260), .B2(new_n1258), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1264), .B(new_n1310), .C1(new_n1266), .C2(new_n1271), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT62), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1305), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1303), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n1272), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1309), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1307), .A2(new_n1317), .ZN(G405));
  AOI21_X1  g1118(.A(G378), .B1(new_n1190), .B2(new_n1220), .ZN(new_n1319));
  OR3_X1    g1119(.A1(new_n1319), .A2(new_n1295), .A3(new_n1289), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1289), .B1(new_n1319), .B2(new_n1295), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1262), .B(new_n1322), .ZN(G402));
endmodule


