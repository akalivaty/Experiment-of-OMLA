//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n204), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(new_n207), .A2(G274), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT69), .B(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G238), .ZN(new_n255));
  INV_X1    g0055(.A(new_n214), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n220), .A2(G1698), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n262), .B1(G226), .B2(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n258), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT13), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n267), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n258), .A2(new_n259), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n253), .B1(new_n270), .B2(G238), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n268), .A2(new_n273), .A3(KEYINPUT72), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT72), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n269), .A2(new_n271), .A3(new_n275), .A4(new_n272), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G169), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT14), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n274), .A2(new_n279), .A3(G169), .A4(new_n276), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n268), .A2(new_n273), .A3(G179), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n208), .A2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n214), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n284), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n214), .A3(new_n289), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n207), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n292), .A2(new_n296), .A3(new_n297), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n282), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n268), .A2(G190), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n304), .B2(new_n273), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n274), .A2(G200), .A3(new_n276), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT7), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n310), .B1(new_n313), .B2(G20), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n263), .A2(new_n264), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n284), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n219), .A2(new_n284), .ZN(new_n318));
  OAI21_X1  g0118(.A(G20), .B1(new_n318), .B2(new_n203), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n283), .A2(G159), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n309), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT7), .B1(new_n315), .B2(new_n208), .ZN(new_n323));
  NOR4_X1   g0123(.A1(new_n263), .A2(new_n264), .A3(new_n310), .A4(G20), .ZN(new_n324));
  OAI21_X1  g0124(.A(G68), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n321), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(KEYINPUT16), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n290), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G1698), .ZN(new_n329));
  OAI211_X1 g0129(.A(G223), .B(new_n329), .C1(new_n263), .C2(new_n264), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT74), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n313), .A2(KEYINPUT74), .A3(G223), .A4(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n329), .B1(new_n311), .B2(new_n312), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n335), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n258), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n254), .B1(new_n220), .B2(new_n260), .ZN(new_n338));
  OAI21_X1  g0138(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n294), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT8), .B(G58), .Z(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n300), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n343), .B2(new_n298), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT73), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT73), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n341), .C1(new_n343), .C2(new_n298), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n253), .B1(new_n270), .B2(G232), .ZN(new_n349));
  OAI211_X1 g0149(.A(G226), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n350));
  INV_X1    g0150(.A(G33), .ZN(new_n351));
  INV_X1    g0151(.A(G87), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n332), .B2(new_n333), .ZN(new_n354));
  OAI211_X1 g0154(.A(G190), .B(new_n349), .C1(new_n354), .C2(new_n258), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n328), .A2(new_n339), .A3(new_n348), .A4(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT17), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n328), .A2(new_n348), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n349), .C1(new_n354), .C2(new_n258), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n337), .A2(new_n338), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n358), .B(new_n360), .C1(G169), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT18), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n345), .A2(new_n347), .ZN(new_n364));
  INV_X1    g0164(.A(new_n290), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n325), .A2(new_n326), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n309), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n367), .B2(new_n327), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n360), .B1(new_n361), .B2(G169), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n357), .A2(new_n363), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n335), .A2(G238), .ZN(new_n374));
  AOI21_X1  g0174(.A(G1698), .B1(new_n311), .B2(new_n312), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G232), .ZN(new_n376));
  INV_X1    g0176(.A(G107), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n374), .B(new_n376), .C1(new_n377), .C2(new_n313), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n253), .B1(new_n270), .B2(G244), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G190), .ZN(new_n387));
  INV_X1    g0187(.A(new_n283), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n340), .A2(new_n388), .B1(new_n208), .B2(new_n286), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n287), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n290), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n286), .B1(new_n207), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n299), .A2(new_n393), .B1(new_n286), .B2(new_n294), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n387), .B(new_n396), .C1(new_n397), .C2(new_n386), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT70), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n375), .A2(new_n399), .A3(G222), .ZN(new_n400));
  OAI211_X1 g0200(.A(G222), .B(new_n329), .C1(new_n263), .C2(new_n264), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT70), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n335), .A2(G223), .B1(new_n315), .B2(G77), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n258), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n253), .B1(new_n270), .B2(G226), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n359), .ZN(new_n409));
  INV_X1    g0209(.A(G150), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n340), .A2(new_n287), .B1(new_n410), .B2(new_n388), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n208), .B1(new_n201), .B2(new_n203), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n290), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G50), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n207), .B2(G20), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n299), .A2(new_n415), .B1(new_n414), .B2(new_n294), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n409), .B(new_n417), .C1(G169), .C2(new_n408), .ZN(new_n418));
  INV_X1    g0218(.A(new_n385), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n384), .B1(new_n380), .B2(new_n381), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n359), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G169), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n383), .A2(new_n422), .A3(new_n385), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n423), .A3(new_n395), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n398), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n403), .A2(new_n404), .ZN(new_n426));
  OAI211_X1 g0226(.A(G190), .B(new_n406), .C1(new_n426), .C2(new_n258), .ZN(new_n427));
  OAI21_X1  g0227(.A(G200), .B1(new_n405), .B2(new_n407), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT9), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n417), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n413), .A2(KEYINPUT9), .A3(new_n416), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n427), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT10), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n430), .A2(new_n431), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT10), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n427), .A4(new_n428), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n308), .A2(new_n373), .A3(new_n425), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT75), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT5), .B(G41), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n441), .A2(new_n443), .B1(new_n256), .B2(new_n257), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n444), .B2(G257), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(new_n440), .A3(G257), .A4(new_n258), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(G274), .A3(new_n443), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT76), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n258), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT75), .B1(new_n453), .B2(new_n222), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT76), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(new_n450), .A4(new_n449), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  OAI211_X1 g0258(.A(G250), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(new_n329), .C1(new_n263), .C2(new_n264), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT4), .B1(new_n375), .B2(G244), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n379), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n359), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n451), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n466), .A3(new_n454), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468));
  AND2_X1   g0268(.A1(G97), .A2(G107), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n377), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n283), .A2(G77), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n377), .B1(new_n314), .B2(new_n316), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n290), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n293), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n207), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n293), .A2(new_n480), .A3(new_n214), .A4(new_n289), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(G97), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n467), .A2(new_n422), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n465), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n483), .ZN(new_n486));
  OAI21_X1  g0286(.A(G107), .B1(new_n323), .B2(new_n324), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n473), .A2(G20), .B1(G77), .B2(new_n283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n489), .B2(new_n290), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n464), .A2(new_n466), .A3(G190), .A4(new_n454), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT77), .ZN(new_n493));
  INV_X1    g0293(.A(new_n464), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n452), .B2(new_n456), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n492), .B(new_n493), .C1(new_n397), .C2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n397), .B1(new_n457), .B2(new_n464), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(new_n491), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT77), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n485), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n289), .A2(new_n214), .B1(G20), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n458), .B(new_n208), .C1(G33), .C2(new_n221), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(KEYINPUT20), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT20), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n294), .A2(new_n501), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n481), .B2(new_n501), .ZN(new_n509));
  OAI21_X1  g0309(.A(G169), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n448), .A2(G270), .A3(new_n258), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n450), .ZN(new_n512));
  OAI211_X1 g0312(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(new_n329), .C1(new_n263), .C2(new_n264), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n313), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n379), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT81), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT81), .B(KEYINPUT21), .C1(new_n510), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n512), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(new_n379), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(G179), .ZN(new_n525));
  INV_X1    g0325(.A(new_n506), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n509), .B1(new_n526), .B2(new_n504), .ZN(new_n527));
  OR3_X1    g0327(.A1(new_n525), .A2(KEYINPUT80), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT80), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n523), .A2(new_n524), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  INV_X1    g0332(.A(G190), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n527), .C1(new_n533), .C2(new_n531), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n522), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G250), .B1(new_n442), .B2(G1), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n379), .A2(new_n537), .B1(new_n442), .B2(new_n250), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n255), .A2(G1698), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n263), .B2(new_n264), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  OAI211_X1 g0342(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT78), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n539), .B(new_n544), .C1(new_n264), .C2(new_n263), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n538), .B1(new_n546), .B2(new_n379), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(KEYINPUT79), .A3(G190), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n379), .ZN(new_n549));
  INV_X1    g0349(.A(new_n538), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(G190), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n547), .A2(new_n397), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n208), .B1(new_n266), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n470), .A2(new_n352), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n208), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n556), .B1(new_n287), .B2(new_n221), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n290), .B1(new_n294), .B2(new_n390), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n482), .A2(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n547), .A2(G169), .ZN(new_n568));
  AOI211_X1 g0368(.A(G179), .B(new_n538), .C1(new_n546), .C2(new_n379), .ZN(new_n569));
  INV_X1    g0369(.A(new_n390), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n482), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n208), .A2(KEYINPUT82), .A3(G87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n315), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n577), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n313), .A2(new_n579), .A3(KEYINPUT22), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n208), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n377), .A2(KEYINPUT23), .A3(G20), .ZN(new_n583));
  INV_X1    g0383(.A(new_n542), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n208), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n578), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(new_n580), .A3(new_n588), .A4(new_n585), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n290), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n377), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n293), .B2(G107), .ZN(new_n594));
  AOI22_X1  g0394(.A1(G107), .A2(new_n482), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n597));
  OAI211_X1 g0397(.A(G250), .B(new_n329), .C1(new_n263), .C2(new_n264), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n379), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n444), .A2(G264), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n450), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n422), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n600), .A2(new_n379), .B1(new_n444), .B2(G264), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n359), .A3(new_n450), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n596), .A2(KEYINPUT83), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(G200), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(G190), .A3(new_n450), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n591), .A2(new_n595), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n365), .B1(new_n587), .B2(new_n589), .ZN(new_n611));
  INV_X1    g0411(.A(new_n595), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n604), .B(new_n606), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n575), .A2(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n439), .A2(new_n500), .A3(new_n536), .A4(new_n617), .ZN(G372));
  AOI21_X1  g0418(.A(KEYINPUT87), .B1(new_n433), .B2(new_n436), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n363), .A2(new_n372), .A3(KEYINPUT86), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT86), .B1(new_n363), .B2(new_n372), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n357), .ZN(new_n627));
  INV_X1    g0427(.A(new_n424), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n307), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n627), .B1(new_n303), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n622), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n418), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n439), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n563), .A2(new_n635), .A3(new_n564), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n563), .B2(new_n564), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n573), .B1(new_n555), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n485), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n551), .B(new_n552), .C1(new_n397), .C2(new_n547), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n565), .B1(new_n643), .B2(new_n548), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n465), .A2(new_n484), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n644), .A2(new_n645), .A3(new_n573), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n642), .B(new_n574), .C1(new_n646), .C2(new_n641), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n638), .B1(new_n643), .B2(new_n548), .ZN(new_n648));
  INV_X1    g0448(.A(new_n610), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n649), .A3(new_n573), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n520), .A2(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n613), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n500), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT85), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n500), .A2(new_n650), .A3(new_n652), .A4(KEYINPUT85), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n633), .B1(new_n634), .B2(new_n657), .ZN(G369));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n535), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n651), .A2(KEYINPUT89), .A3(new_n534), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n527), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n660), .A2(new_n661), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT88), .B1(new_n651), .B2(new_n670), .ZN(new_n672));
  OR3_X1    g0472(.A1(new_n651), .A2(KEYINPUT88), .A3(new_n670), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n668), .B1(new_n591), .B2(new_n595), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n616), .A2(new_n675), .B1(new_n613), .B2(new_n668), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(G330), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT90), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n674), .A2(KEYINPUT90), .A3(G330), .A4(new_n676), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n522), .A2(new_n530), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n668), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n683), .A2(new_n616), .B1(new_n613), .B2(new_n667), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n681), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n211), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n558), .A2(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n217), .B2(new_n688), .ZN(new_n691));
  XOR2_X1   g0491(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n692));
  XNOR2_X1  g0492(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G330), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n517), .A2(new_n547), .A3(G179), .A4(new_n605), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n467), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n547), .A2(new_n605), .ZN(new_n698));
  INV_X1    g0498(.A(new_n467), .ZN(new_n699));
  INV_X1    g0499(.A(new_n525), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT30), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n547), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n359), .A3(new_n531), .A4(new_n603), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n697), .B(new_n701), .C1(new_n495), .C2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT31), .B1(new_n704), .B2(new_n667), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n704), .A2(new_n667), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT92), .B(KEYINPUT31), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n617), .A2(new_n500), .A3(new_n536), .A4(new_n668), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n694), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n713), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n485), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n640), .A2(KEYINPUT26), .A3(new_n485), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n522), .A2(new_n607), .A3(new_n530), .A4(new_n615), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n500), .A2(new_n650), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n574), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n668), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n719), .A2(new_n574), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n640), .A2(new_n713), .A3(KEYINPUT26), .A4(new_n485), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n567), .A2(new_n485), .A3(new_n574), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT93), .B1(new_n726), .B2(new_n641), .ZN(new_n727));
  INV_X1    g0527(.A(new_n716), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT94), .A3(new_n668), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n712), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n657), .A2(new_n667), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n711), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n693), .B1(new_n736), .B2(G1), .ZN(G364));
  AND2_X1   g0537(.A1(new_n674), .A2(G330), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n208), .A2(G13), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n207), .B1(new_n739), .B2(G45), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n688), .A2(KEYINPUT95), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  INV_X1    g0542(.A(new_n740), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n687), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n674), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n214), .B1(G20), .B2(new_n422), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n208), .A2(new_n359), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n533), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT98), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G326), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(G190), .A3(new_n397), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n756), .A2(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n208), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n758), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n313), .B(new_n761), .C1(G329), .C2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n533), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n208), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n768), .A2(G294), .B1(new_n770), .B2(G303), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n752), .A2(G190), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n762), .A2(new_n533), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n772), .A2(new_n773), .B1(new_n775), .B2(G283), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n755), .A2(new_n765), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n753), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n778), .A2(new_n414), .B1(new_n774), .B2(new_n377), .ZN(new_n779));
  INV_X1    g0579(.A(new_n772), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n780), .A2(new_n284), .B1(new_n769), .B2(new_n352), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n767), .B(KEYINPUT97), .Z(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G97), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n763), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n313), .B1(new_n756), .B2(new_n219), .ZN(new_n788));
  INV_X1    g0588(.A(new_n759), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G77), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n782), .A2(new_n784), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n750), .B1(new_n777), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n686), .A2(new_n315), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(G355), .B1(new_n501), .B2(new_n686), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n248), .A2(G45), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n686), .A2(new_n313), .ZN(new_n796));
  INV_X1    g0596(.A(new_n251), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n217), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT96), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n749), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n799), .B2(KEYINPUT96), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n792), .B(new_n745), .C1(new_n800), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n803), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n674), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n748), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n424), .A2(KEYINPUT101), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT101), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n421), .A2(new_n423), .A3(new_n813), .A4(new_n395), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n395), .A2(new_n667), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT102), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n398), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n628), .A2(new_n667), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR3_X1    g0619(.A1(new_n733), .A2(KEYINPUT103), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT103), .B1(new_n733), .B2(new_n819), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n657), .A2(new_n667), .A3(new_n817), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n746), .B1(new_n823), .B2(new_n711), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n711), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n749), .A2(new_n801), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n746), .B1(G77), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT100), .ZN(new_n829));
  INV_X1    g0629(.A(new_n756), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(G143), .B1(new_n789), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n778), .B2(new_n832), .C1(new_n410), .C2(new_n780), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n774), .A2(new_n284), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n315), .B(new_n837), .C1(G132), .C2(new_n764), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n768), .A2(G58), .B1(new_n770), .B2(G50), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n756), .A2(new_n841), .B1(new_n759), .B2(new_n501), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n313), .B(new_n842), .C1(G311), .C2(new_n764), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n772), .A2(G283), .B1(new_n753), .B2(G303), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n774), .A2(new_n352), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G107), .B2(new_n770), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n784), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n829), .B1(new_n750), .B2(new_n848), .C1(new_n819), .C2(new_n802), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n825), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  NAND2_X1  g0651(.A1(new_n302), .A2(new_n667), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n303), .A2(new_n307), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n307), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n302), .B(new_n667), .C1(new_n854), .C2(new_n282), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n853), .A2(new_n855), .B1(new_n817), .B2(new_n818), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n707), .B1(new_n704), .B2(new_n667), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(KEYINPUT31), .B2(new_n706), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n709), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT106), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n665), .B1(new_n328), .B2(new_n348), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(KEYINPUT104), .B(new_n665), .C1(new_n328), .C2(new_n348), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n356), .B(new_n362), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n665), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n358), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n356), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n370), .A2(KEYINPUT37), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n866), .A2(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT104), .B1(new_n368), .B2(new_n665), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n862), .A2(new_n863), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n872), .A2(new_n873), .B1(new_n373), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n356), .B1(new_n368), .B2(new_n369), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n869), .A2(new_n370), .A3(KEYINPUT37), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT105), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n373), .A2(new_n877), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n870), .A2(new_n871), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n880), .B1(new_n874), .B2(new_n875), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n887), .B(new_n873), .C1(new_n888), .C2(new_n879), .ZN(new_n889));
  AND4_X1   g0689(.A1(KEYINPUT38), .A2(new_n884), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n861), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n884), .A2(new_n886), .A3(new_n889), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT38), .A4(new_n886), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n860), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(KEYINPUT40), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT86), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n869), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n362), .A2(new_n356), .A3(new_n868), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n870), .A2(new_n899), .A3(KEYINPUT37), .A4(new_n362), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n362), .A2(KEYINPUT18), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n370), .A2(new_n371), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n363), .A2(new_n372), .A3(KEYINPUT86), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n357), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n904), .B1(new_n909), .B2(new_n862), .ZN(new_n910));
  XOR2_X1   g0710(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n895), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n898), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n439), .A2(new_n859), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n917), .A2(new_n918), .A3(new_n694), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n891), .A2(new_n896), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n853), .A2(new_n855), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n812), .A2(new_n814), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n668), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n822), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n868), .B1(new_n625), .B2(new_n357), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n911), .B1(new_n926), .B2(new_n904), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT108), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n895), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n303), .A2(new_n667), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n895), .C1(new_n910), .C2(new_n912), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n929), .B1(new_n894), .B2(new_n895), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n930), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n626), .A2(new_n665), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n925), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n732), .A2(new_n734), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n632), .B1(new_n938), .B2(new_n439), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n919), .A2(new_n940), .B1(new_n207), .B2(new_n739), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n919), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n501), .B(new_n216), .C1(new_n473), .C2(KEYINPUT35), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(KEYINPUT35), .B2(new_n473), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT36), .Z(new_n945));
  OR3_X1    g0745(.A1(new_n217), .A2(new_n286), .A3(new_n318), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n201), .A2(G68), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n207), .B(G13), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n942), .A2(new_n945), .A3(new_n948), .ZN(G367));
  INV_X1    g0749(.A(KEYINPUT109), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n490), .A2(new_n668), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n500), .A2(new_n951), .B1(new_n485), .B2(new_n667), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n684), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n684), .A2(new_n952), .A3(new_n950), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n684), .A2(new_n952), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n684), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n684), .A2(new_n952), .A3(new_n950), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n953), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n956), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n679), .A2(KEYINPUT110), .A3(new_n680), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n676), .B1(new_n682), .B2(new_n668), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n683), .A2(new_n616), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n738), .B(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n736), .A3(KEYINPUT111), .A4(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT111), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n681), .A2(new_n964), .A3(KEYINPUT110), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n965), .A2(new_n963), .A3(new_n960), .A4(new_n956), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n970), .B(new_n711), .C1(new_n732), .C2(new_n734), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n735), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n687), .B(KEYINPUT41), .Z(new_n979));
  OAI21_X1  g0779(.A(new_n740), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n496), .A2(new_n499), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n607), .A2(new_n615), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n667), .B1(new_n983), .B2(new_n645), .ZN(new_n984));
  INV_X1    g0784(.A(new_n952), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n968), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n984), .B1(new_n986), .B2(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT42), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n638), .A2(new_n667), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n574), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n640), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n988), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n989), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n681), .A2(new_n985), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n980), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n796), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n804), .B1(new_n211), .B2(new_n390), .C1(new_n999), .C2(new_n238), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n754), .A2(G143), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT114), .B(G137), .Z(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n763), .B1(new_n759), .B2(new_n201), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n315), .B(new_n1003), .C1(G150), .C2(new_n830), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n769), .A2(new_n219), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n774), .A2(new_n286), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G159), .C2(new_n772), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n783), .A2(G68), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1001), .A2(new_n1004), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT113), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT112), .B(G317), .Z(new_n1011));
  OAI221_X1 g0811(.A(new_n315), .B1(new_n774), .B2(new_n221), .C1(new_n763), .C2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n754), .A2(G311), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n770), .A2(G116), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT46), .ZN(new_n1016));
  INV_X1    g0816(.A(G283), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n756), .A2(new_n515), .B1(new_n759), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G107), .B2(new_n768), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(new_n841), .C2(new_n780), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1009), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT47), .Z(new_n1022));
  OAI211_X1 g0822(.A(new_n746), .B(new_n1000), .C1(new_n1022), .C2(new_n750), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n992), .A2(new_n803), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n998), .A2(new_n1026), .ZN(G387));
  OR2_X1    g0827(.A1(new_n676), .A2(new_n808), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n796), .B1(new_n235), .B2(new_n251), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n793), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n689), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n340), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g0833(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n689), .A3(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1031), .A2(new_n1035), .B1(new_n377), .B2(new_n686), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n746), .B1(new_n1036), .B2(new_n805), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT115), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n756), .A2(new_n414), .B1(new_n759), .B2(new_n284), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n315), .B(new_n1039), .C1(G150), .C2(new_n764), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n783), .A2(new_n570), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n753), .A2(G159), .B1(new_n775), .B2(G97), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n772), .A2(new_n342), .B1(new_n770), .B2(G77), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(KEYINPUT116), .B(G322), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n754), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1011), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n830), .A2(new_n1047), .B1(new_n789), .B2(G303), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(new_n760), .C2(new_n780), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n767), .A2(new_n1017), .B1(new_n769), .B2(new_n841), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(KEYINPUT49), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n313), .B1(new_n764), .B2(G326), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n501), .C2(new_n774), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT49), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1044), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1038), .B1(new_n749), .B2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n970), .A2(new_n743), .B1(new_n1028), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n736), .A2(new_n970), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n976), .A2(new_n687), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n243), .A2(new_n796), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n805), .B1(G97), .B2(new_n686), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n745), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n315), .B(new_n845), .C1(new_n342), .C2(new_n789), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n770), .A2(G68), .B1(new_n764), .B2(G143), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1067), .B1(KEYINPUT118), .B2(new_n1069), .C1(new_n201), .C2(new_n780), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n753), .B1(new_n830), .B2(G159), .ZN(new_n1071));
  XOR2_X1   g0871(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1069), .A2(KEYINPUT118), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n783), .A2(G77), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n313), .B1(new_n764), .B2(new_n1045), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n377), .B2(new_n774), .C1(new_n1017), .C2(new_n769), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT119), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n767), .A2(new_n501), .B1(new_n759), .B2(new_n841), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G317), .A2(new_n753), .B1(new_n830), .B2(G311), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(G303), .C2(new_n772), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1078), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1066), .B1(new_n750), .B2(new_n1086), .C1(new_n985), .C2(new_n808), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n681), .B(new_n964), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n740), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n971), .A2(new_n977), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n688), .B1(new_n1088), .B2(new_n976), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G390));
  INV_X1    g0893(.A(new_n931), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n913), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT94), .B1(new_n730), .B2(new_n668), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n722), .B(new_n667), .C1(new_n724), .C2(new_n729), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n819), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n923), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1095), .B1(new_n1099), .B2(new_n921), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT39), .B1(new_n885), .B2(new_n890), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(KEYINPUT108), .A3(new_n932), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n657), .A2(new_n667), .A3(new_n817), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n923), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n921), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1102), .A2(new_n930), .B1(new_n1105), .B2(new_n1094), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n708), .A2(new_n709), .ZN(new_n1107));
  AND4_X1   g0907(.A1(G330), .A2(new_n1107), .A3(new_n819), .A4(new_n921), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1100), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n694), .B1(new_n858), .B2(new_n709), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n856), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1095), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n723), .A2(new_n731), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1104), .B1(new_n1113), .B2(new_n819), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n921), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1105), .A2(new_n1094), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1111), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n710), .A2(new_n819), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1111), .B1(new_n1121), .B2(new_n921), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n924), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n921), .B1(new_n1110), .B2(new_n819), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1108), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1098), .A2(new_n923), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT120), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1098), .A2(new_n1126), .A3(new_n1129), .A4(new_n923), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1124), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1113), .A2(KEYINPUT29), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n734), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n439), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n439), .A2(new_n1110), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n633), .A3(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1109), .A2(new_n1120), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1123), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1111), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1108), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1116), .A2(new_n1119), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1136), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1137), .A2(new_n1145), .A3(new_n687), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1141), .A2(new_n743), .A3(new_n1143), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1117), .A2(new_n801), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n746), .B1(new_n342), .B2(new_n827), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT121), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n759), .A2(new_n221), .B1(new_n763), .B2(new_n841), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n313), .B(new_n1151), .C1(G116), .C2(new_n830), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n837), .B1(G87), .B2(new_n770), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n772), .A2(G107), .B1(new_n753), .B2(G283), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1152), .A2(new_n1076), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n769), .A2(new_n410), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n315), .B1(new_n775), .B2(new_n202), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n783), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1157), .B1(KEYINPUT122), .B2(new_n1158), .C1(new_n1159), .C2(new_n785), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1002), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1162), .A2(new_n772), .B1(new_n753), .B2(G128), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n830), .A2(G132), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT54), .B(G143), .Z(new_n1165));
  AOI22_X1  g0965(.A1(new_n789), .A2(new_n1165), .B1(new_n764), .B2(G125), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1155), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1150), .B1(new_n749), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1148), .A2(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1147), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1146), .A2(new_n1171), .ZN(G378));
  OAI21_X1  g0972(.A(new_n746), .B1(new_n202), .B2(new_n827), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n417), .A2(new_n867), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n622), .B2(new_n418), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT87), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n418), .B(new_n1176), .C1(new_n1178), .C2(new_n619), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1175), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n418), .B1(new_n1178), .B2(new_n619), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n417), .A3(new_n867), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1179), .A3(new_n1174), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1181), .A2(KEYINPUT123), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT123), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1187), .A2(new_n802), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n414), .B1(G33), .B2(G41), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n315), .B2(new_n252), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n221), .A2(new_n780), .B1(new_n778), .B2(new_n501), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n219), .A2(new_n774), .B1(new_n769), .B2(new_n286), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G41), .B(new_n313), .C1(new_n764), .C2(G283), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n830), .A2(G107), .B1(new_n789), .B2(new_n570), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1193), .A2(new_n1008), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT58), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1190), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n756), .A2(new_n1199), .B1(new_n759), .B2(new_n832), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G132), .B2(new_n772), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n753), .A2(G125), .B1(new_n770), .B2(new_n1165), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n1159), .C2(new_n410), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n775), .A2(G159), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1198), .B1(new_n1197), .B2(new_n1196), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1173), .B(new_n1188), .C1(new_n749), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n913), .A2(new_n914), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(G330), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1187), .B(new_n1213), .C1(new_n897), .C2(KEYINPUT40), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n860), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n896), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT106), .B1(new_n894), .B2(new_n895), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT40), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1212), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1181), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1184), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1214), .B(new_n937), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1223), .B1(new_n898), .B2(new_n1212), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n937), .B1(new_n1227), .B2(new_n1214), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1210), .B1(new_n1229), .B2(new_n743), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1109), .A2(new_n1120), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1136), .B1(new_n1231), .B2(new_n1139), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n937), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1214), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n687), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1144), .B1(new_n1239), .B2(new_n1131), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1229), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1230), .B1(new_n1238), .B2(new_n1241), .ZN(G375));
  NAND2_X1  g1042(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n979), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1115), .A2(new_n801), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n746), .B1(G68), .B2(new_n827), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n756), .A2(new_n1017), .B1(new_n759), .B2(new_n377), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n313), .B(new_n1249), .C1(G303), .C2(new_n764), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1006), .B1(G116), .B2(new_n772), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n753), .A2(G294), .B1(new_n770), .B2(G97), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1041), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n772), .A2(new_n1165), .B1(new_n775), .B2(G58), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n785), .B2(new_n769), .C1(new_n1159), .C2(new_n414), .ZN(new_n1255));
  INV_X1    g1055(.A(G132), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n778), .A2(KEYINPUT124), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT124), .B1(new_n778), .B2(new_n1256), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n315), .B1(new_n789), .B2(G150), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n830), .A2(new_n1162), .B1(new_n764), .B2(G128), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1253), .B1(new_n1255), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1248), .B1(new_n1262), .B2(new_n749), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1247), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1131), .B2(new_n740), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(new_n1266), .ZN(G381));
  OR4_X1    g1067(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1268), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1269));
  INV_X1    g1069(.A(G375), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G407));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n666), .A2(G213), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G375), .C2(new_n1275), .ZN(G409));
  OAI211_X1 g1076(.A(G378), .B(new_n1230), .C1(new_n1238), .C2(new_n1241), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1240), .A2(new_n1229), .A3(new_n1244), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1230), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1272), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1274), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n1136), .A4(new_n1123), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n687), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT60), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1245), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1288), .B2(new_n1266), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1265), .B(new_n850), .C1(new_n1285), .C2(new_n1287), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1282), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1284), .B1(new_n1245), .B2(new_n1286), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n850), .B1(new_n1292), .B2(new_n1265), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1288), .A2(G384), .A3(new_n1266), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(KEYINPUT125), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1281), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1274), .A2(G2897), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1293), .A2(KEYINPUT125), .A3(new_n1294), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT125), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1273), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1299), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1302), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1281), .A2(new_n1296), .A3(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1298), .A2(new_n1307), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G390), .B1(new_n998), .B2(new_n1026), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n1025), .B(new_n1092), .C1(new_n980), .C2(new_n997), .ZN(new_n1313));
  OAI21_X1  g1113(.A(KEYINPUT126), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(new_n810), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  OAI211_X1 g1117(.A(KEYINPUT126), .B(new_n1317), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1316), .A2(new_n1318), .A3(KEYINPUT127), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT127), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1281), .A2(new_n1305), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1302), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1297), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1281), .A2(new_n1296), .A3(KEYINPUT63), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1324), .A2(new_n1325), .A3(new_n1327), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1322), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1272), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1277), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1296), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1331), .B(new_n1277), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1321), .A2(new_n1335), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1333), .B(new_n1334), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(G402));
endmodule


