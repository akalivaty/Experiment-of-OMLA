//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n451, new_n453,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n450));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  INV_X1    g027(.A(new_n451), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n453), .A2(G567), .ZN(G234));
  NAND2_X1  g029(.A1(new_n453), .A2(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XOR2_X1   g031(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n457));
  XNOR2_X1  g032(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  NAND2_X1  g037(.A1(new_n458), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G567), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(KEYINPUT3), .A3(new_n477), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n481), .A2(G137), .A3(new_n482), .A4(new_n468), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n481), .A2(new_n468), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n486), .A2(new_n482), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n482), .A2(G138), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n481), .A2(new_n468), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n468), .A2(new_n470), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n482), .A3(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n481), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n506), .B(G2104), .C1(G114), .C2(new_n482), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n495), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n502), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n507), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT71), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT5), .B1(new_n515), .B2(KEYINPUT72), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT73), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G62), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G88), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G50), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR3_X1    g104(.A1(new_n523), .A2(new_n529), .A3(KEYINPUT75), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT75), .B1(new_n523), .B2(new_n529), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(KEYINPUT76), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n534), .A2(G543), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n519), .A2(new_n520), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n525), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n519), .A2(new_n520), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n546), .A2(G63), .A3(G651), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n540), .A2(new_n543), .A3(new_n545), .A4(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n524), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n538), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n546), .A2(G64), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n514), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n539), .A2(G43), .B1(new_n542), .B2(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n541), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND4_X1  g144(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n537), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n541), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n542), .B2(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n542), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n546), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n538), .ZN(G288));
  NAND3_X1  g157(.A1(new_n519), .A2(G61), .A3(new_n520), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n514), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n519), .A2(G86), .A3(new_n520), .ZN(new_n586));
  NAND2_X1  g161(.A1(G48), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n525), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n539), .A2(G47), .B1(new_n542), .B2(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n546), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n514), .B2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n542), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n541), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(G54), .A2(new_n539), .B1(new_n600), .B2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n594), .B1(new_n603), .B2(G868), .ZN(G321));
  XOR2_X1   g179(.A(G321), .B(KEYINPUT77), .Z(G284));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  XOR2_X1   g184(.A(KEYINPUT78), .B(G559), .Z(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(G860), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT79), .ZN(G148));
  NOR2_X1   g187(.A1(new_n563), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n603), .A2(new_n610), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n613), .B1(new_n616), .B2(G868), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g194(.A1(new_n478), .A2(new_n468), .A3(new_n470), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT82), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n487), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n489), .A2(G123), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  OAI22_X1  g205(.A1(new_n622), .A2(new_n623), .B1(G2096), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G2096), .B2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT84), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(KEYINPUT14), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT86), .Z(new_n657));
  NOR2_X1   g232(.A1(G2072), .A2(G2078), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n444), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(KEYINPUT17), .Z(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n662), .B2(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n656), .A3(new_n655), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n657), .A3(new_n655), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n623), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT87), .B(G2096), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OR3_X1    g252(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT89), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n671), .A3(new_n672), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n671), .B(new_n672), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n681), .B(new_n682), .C1(new_n677), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G23), .ZN(new_n692));
  INV_X1    g267(.A(G288), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT33), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n691), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G1971), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT32), .B(G1981), .ZN(new_n701));
  NOR2_X1   g276(.A1(G6), .A2(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n589), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT93), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n704), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n696), .B(new_n705), .C1(new_n701), .C2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT34), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  OR2_X1    g284(.A1(G25), .A2(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n487), .A2(G131), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n482), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n489), .A2(G119), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n710), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n691), .A2(G24), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT92), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G290), .B2(G16), .ZN(new_n725));
  INV_X1    g300(.A(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n720), .A2(new_n721), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n708), .A2(new_n709), .A3(new_n722), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n719), .A2(G33), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n487), .A2(G139), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G127), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n499), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT98), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n482), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n733), .B1(new_n744), .B2(new_n719), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT99), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n719), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n719), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT101), .B(G2078), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n719), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n487), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n489), .A2(G128), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n482), .A2(G116), .ZN(new_n757));
  OAI21_X1  g332(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n754), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n747), .A2(new_n751), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n691), .A2(G19), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT95), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n564), .B2(new_n691), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G1341), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n691), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n691), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n719), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n487), .A2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n489), .A2(G129), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(G105), .A2(new_n478), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n775), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n719), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT27), .B(G1996), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT24), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT24), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n484), .B2(new_n719), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT31), .B(G11), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n719), .B1(new_n795), .B2(G28), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(KEYINPUT100), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(G28), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n796), .B2(KEYINPUT100), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n794), .B1(new_n797), .B2(new_n799), .C1(new_n630), .C2(new_n719), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n792), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n769), .A2(new_n773), .A3(new_n786), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT94), .B(G1348), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n603), .A2(G16), .ZN(new_n804));
  OR2_X1    g379(.A1(G4), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n691), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n691), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1966), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n804), .A2(new_n805), .A3(new_n803), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n802), .A2(new_n806), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n691), .A2(G20), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT23), .Z(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G299), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(G1956), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n719), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n719), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT29), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n819), .B2(G2090), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n811), .B(new_n820), .C1(G2090), .C2(new_n819), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n732), .A2(new_n765), .A3(new_n821), .ZN(G311));
  OR3_X1    g397(.A1(new_n732), .A2(new_n765), .A3(new_n821), .ZN(G150));
  NAND2_X1  g398(.A1(new_n603), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n550), .A2(new_n826), .B1(new_n827), .B2(new_n538), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n546), .A2(G67), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n514), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n564), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n563), .B1(new_n831), .B2(new_n828), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n825), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n832), .A2(new_n839), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n718), .B(new_n621), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n744), .B(new_n782), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n504), .A2(new_n508), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n762), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n762), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n487), .A2(G142), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT102), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n489), .A2(G130), .ZN(new_n854));
  OR2_X1    g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G118), .C2(new_n482), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n850), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n850), .B2(new_n851), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n848), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n847), .A2(new_n859), .A3(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n630), .B(new_n484), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n493), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n862), .A2(new_n866), .A3(new_n863), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n835), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n616), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n602), .B(G299), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT41), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n876), .B(KEYINPUT104), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(G166), .B(new_n693), .ZN(new_n882));
  XNOR2_X1  g457(.A(G290), .B(G305), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n878), .B2(new_n880), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n881), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(G868), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g464(.A(new_n888), .B1(G868), .B2(new_n832), .ZN(G331));
  INV_X1    g465(.A(new_n876), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n835), .B(G301), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(G168), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n836), .A2(G301), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n835), .A2(G171), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(G286), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n891), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(G168), .ZN(new_n898));
  OAI21_X1  g473(.A(G286), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n877), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n900), .A3(new_n884), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n869), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n884), .B1(new_n897), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n901), .A2(new_n869), .ZN(new_n905));
  INV_X1    g480(.A(new_n884), .ZN(new_n906));
  INV_X1    g481(.A(new_n900), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n904), .B1(new_n910), .B2(KEYINPUT43), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n897), .A2(new_n900), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n906), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n869), .A4(new_n901), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT105), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n905), .A2(new_n919), .A3(new_n916), .A4(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n912), .B1(new_n910), .B2(KEYINPUT43), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT106), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT106), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(G397));
  NOR2_X1   g500(.A1(G290), .A2(G1986), .ZN(new_n926));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n510), .B2(new_n511), .ZN(new_n928));
  XOR2_X1   g503(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n474), .A2(G40), .A3(new_n483), .A4(new_n479), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT48), .Z(new_n934));
  XOR2_X1   g509(.A(new_n762), .B(G2067), .Z(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n782), .B(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n718), .B(new_n721), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n934), .B1(new_n940), .B2(new_n932), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n936), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT46), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n935), .A2(new_n783), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(new_n932), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n938), .A2(new_n713), .A3(new_n717), .A4(new_n721), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G2067), .B2(new_n762), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n941), .B(new_n946), .C1(new_n932), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT125), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT49), .ZN(new_n951));
  OAI21_X1  g526(.A(G1981), .B1(new_n585), .B2(new_n588), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT110), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n954), .B(G1981), .C1(new_n585), .C2(new_n588), .ZN(new_n955));
  XOR2_X1   g530(.A(KEYINPUT109), .B(G1981), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n589), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n951), .ZN(new_n962));
  OAI21_X1  g537(.A(G8), .B1(new_n928), .B2(new_n931), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT108), .B(G8), .C1(new_n928), .C2(new_n931), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n965), .A2(new_n966), .B1(G1976), .B2(new_n693), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n693), .A2(G1976), .ZN(new_n972));
  INV_X1    g547(.A(G1976), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(G288), .B2(new_n973), .ZN(new_n974));
  AND4_X1   g549(.A1(G40), .A2(new_n474), .A3(new_n483), .A4(new_n479), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n849), .A2(new_n975), .A3(new_n927), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT108), .B1(new_n976), .B2(G8), .ZN(new_n977));
  INV_X1    g552(.A(new_n966), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n972), .B(new_n974), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n968), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n504), .B2(new_n508), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n931), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G2090), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n504), .A2(new_n508), .A3(new_n495), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT71), .B1(new_n510), .B2(new_n511), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n983), .B(new_n984), .C1(new_n987), .C2(new_n982), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n975), .B1(new_n928), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n927), .B1(new_n509), .B2(new_n512), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n929), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n992), .B2(G1971), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(G166), .B2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n530), .A2(KEYINPUT55), .A3(G8), .A4(new_n531), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n998), .A3(G8), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n993), .B2(G8), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n980), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n983), .B(new_n791), .C1(new_n987), .C2(new_n982), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n929), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n987), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n931), .B1(new_n928), .B2(new_n989), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1966), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G286), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(KEYINPUT63), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n958), .A2(new_n959), .A3(new_n951), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n965), .A2(new_n966), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(new_n960), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n979), .B1(new_n970), .B2(new_n969), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT115), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n968), .A2(new_n971), .A3(new_n1017), .A4(new_n979), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n931), .B1(new_n928), .B2(KEYINPUT50), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(KEYINPUT114), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n982), .B(new_n927), .C1(new_n509), .C2(new_n512), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT114), .B(new_n975), .C1(new_n981), .C2(new_n982), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n984), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n931), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n987), .B2(new_n1005), .ZN(new_n1027));
  INV_X1    g602(.A(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n998), .B1(new_n1030), .B2(G8), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n1000), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1019), .A2(new_n1020), .A3(new_n1032), .A4(new_n1010), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n995), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n999), .B1(new_n1036), .B2(new_n998), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1020), .B1(new_n1038), .B2(new_n1010), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1011), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G286), .A2(G8), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1009), .A2(KEYINPUT51), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  AOI211_X1 g619(.A(G1384), .B(new_n929), .C1(new_n985), .C2(new_n986), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1007), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1003), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1043), .B(G8), .C1(new_n1048), .C2(G286), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1041), .B1(new_n1047), .B2(new_n1003), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT123), .B(new_n1041), .C1(new_n1047), .C2(new_n1003), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1042), .B(new_n1049), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1050), .B(new_n1051), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(KEYINPUT62), .A3(new_n1042), .A4(new_n1049), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1027), .B2(G2078), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n983), .B1(new_n987), .B2(new_n982), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n772), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1006), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1007), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G171), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1066), .B(new_n1037), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G288), .A2(G1976), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n968), .A2(new_n1068), .B1(new_n589), .B2(new_n956), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n967), .B(KEYINPUT112), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1069), .A2(new_n1070), .B1(new_n980), .B2(new_n999), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g648(.A(KEYINPUT113), .B1(new_n980), .B2(new_n999), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1059), .A2(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1021), .A2(KEYINPUT114), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n815), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n992), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G299), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n607), .A2(KEYINPUT57), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G299), .A2(KEYINPUT119), .A3(new_n1082), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n975), .B1(new_n928), .B2(KEYINPUT50), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G1348), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n976), .A2(G2067), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT121), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1062), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1090), .B1(new_n1100), .B2(new_n602), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1078), .A2(new_n1088), .A3(new_n1080), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1078), .A2(new_n1088), .A3(KEYINPUT120), .A4(new_n1080), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT121), .B(new_n1094), .C1(new_n1062), .C2(new_n1096), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT60), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n603), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n976), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT58), .B(G1341), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1027), .A2(G1996), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n564), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1121), .A3(new_n564), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1090), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1088), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1123), .B(new_n1124), .C1(new_n1126), .C2(KEYINPUT61), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1115), .B1(new_n1127), .B2(KEYINPUT122), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1130), .A2(new_n1102), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1131), .B(new_n1132), .C1(KEYINPUT61), .C2(new_n1126), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1108), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1065), .A2(G171), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1026), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n930), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1061), .A2(new_n1063), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G171), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(KEYINPUT124), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(KEYINPUT124), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT54), .B(new_n1135), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1066), .B1(G171), .B2(new_n1137), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1141), .A2(new_n1144), .A3(new_n1038), .A4(new_n1054), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1040), .B(new_n1075), .C1(new_n1134), .C2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n938), .A2(new_n939), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G290), .B(new_n726), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n932), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n950), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT61), .B1(new_n1106), .B2(new_n1090), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1124), .A2(new_n1123), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT122), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1115), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1133), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1145), .B1(new_n1156), .B2(new_n1107), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1040), .A2(new_n1075), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n950), .B(new_n1150), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n949), .B1(new_n1151), .B2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g736(.A1(G227), .A2(new_n465), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n653), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g738(.A1(G229), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g739(.A1(new_n1165), .A2(new_n871), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n911), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g741(.A(new_n1167), .B(KEYINPUT126), .ZN(G308));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1169));
  XNOR2_X1  g743(.A(new_n1167), .B(new_n1169), .ZN(G225));
endmodule


