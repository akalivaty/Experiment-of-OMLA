//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(KEYINPUT76), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT76), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G155gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n208), .B1(new_n220), .B2(G162gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n207), .A2(new_n212), .A3(new_n214), .A4(new_n209), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n204), .B(new_n216), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT77), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT76), .B(G155gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n225), .B2(new_n211), .ZN(new_n226));
  INV_X1    g025(.A(new_n222), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n228), .A2(new_n229), .A3(new_n204), .A4(new_n216), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G134gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n237), .B(new_n240), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244));
  INV_X1    g043(.A(G120gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G113gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT1), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n236), .B(KEYINPUT68), .C1(new_n238), .C2(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n243), .A2(new_n251), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n203), .B1(new_n231), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n226), .A2(new_n227), .B1(new_n215), .B2(new_n210), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n251), .A3(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n255), .A2(new_n251), .A3(new_n243), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT5), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n251), .A2(new_n243), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n252), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n256), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(new_n203), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(KEYINPUT78), .A3(new_n259), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n259), .A2(KEYINPUT78), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n272), .A3(new_n262), .A4(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n271), .B1(new_n267), .B2(new_n274), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI211_X1 g078(.A(new_n276), .B(new_n271), .C1(new_n267), .C2(new_n274), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT26), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(KEYINPUT28), .A3(new_n293), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n290), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n307), .A2(new_n308), .B1(new_n310), .B2(new_n293), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT25), .B1(new_n313), .B2(G169gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n288), .B1(KEYINPUT23), .B2(new_n286), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n290), .A2(new_n304), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n293), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n307), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n282), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n284), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n320), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n317), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n317), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n299), .B(new_n301), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n301), .A2(KEYINPUT29), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n312), .A2(new_n316), .B1(new_n329), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n298), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G218gat), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT72), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT72), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G197gat), .B(G204gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G211gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n340), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n347), .B1(new_n351), .B2(KEYINPUT22), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT22), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT71), .B(G211gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n340), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n341), .A2(new_n343), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n347), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n337), .A2(new_n298), .A3(new_n300), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n334), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n337), .A2(new_n332), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n298), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(new_n301), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n361), .B(new_n363), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT83), .B(KEYINPUT37), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n360), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(KEYINPUT38), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n339), .A2(new_n361), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n359), .B(new_n363), .C1(new_n366), .C2(new_n370), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT37), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT82), .A4(KEYINPUT37), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n360), .A2(new_n371), .A3(new_n376), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(new_n360), .B2(new_n371), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT38), .B1(new_n378), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n281), .A2(new_n387), .A3(new_n388), .A4(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n360), .A2(new_n371), .A3(KEYINPUT30), .A4(new_n376), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n299), .B1(new_n333), .B2(new_n334), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n359), .B(new_n362), .C1(new_n394), .C2(new_n369), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n361), .B1(new_n335), .B2(new_n338), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n377), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT74), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n393), .B1(new_n397), .B2(KEYINPUT74), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n388), .A2(KEYINPUT75), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT75), .B1(new_n388), .B2(new_n400), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n398), .A2(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT40), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n231), .A2(new_n253), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n272), .A2(new_n273), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT39), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n203), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n271), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT39), .B1(new_n265), .B2(new_n203), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n406), .B2(new_n203), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n411), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n413), .A2(KEYINPUT40), .A3(new_n271), .A4(new_n408), .ZN(new_n414));
  INV_X1    g213(.A(new_n278), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n403), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n231), .A2(new_n367), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n361), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n353), .B2(new_n358), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n204), .B1(new_n421), .B2(KEYINPUT80), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n423), .B(KEYINPUT29), .C1(new_n353), .C2(new_n358), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n252), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G22gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n359), .B1(new_n231), .B2(new_n367), .ZN(new_n428));
  INV_X1    g227(.A(new_n358), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n357), .B1(new_n356), .B2(new_n347), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n367), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n255), .B1(new_n431), .B2(new_n204), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n418), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n427), .B1(new_n426), .B2(new_n433), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n426), .A2(new_n438), .A3(new_n433), .A4(new_n427), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT31), .B(G50gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  XOR2_X1   g242(.A(new_n443), .B(KEYINPUT79), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n436), .A2(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n434), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n392), .A2(new_n417), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n451));
  INV_X1    g250(.A(new_n263), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n394), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G227gat), .ZN(new_n454));
  INV_X1    g253(.A(G233gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n299), .B(new_n263), .C1(new_n333), .C2(new_n334), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(G15gat), .B(G43gat), .Z(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n453), .A2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(new_n456), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n458), .A2(KEYINPUT32), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n463), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n458), .B2(new_n459), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  AOI211_X1 g275(.A(KEYINPUT34), .B(new_n456), .C1(new_n453), .C2(new_n457), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n471), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n471), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n451), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n478), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n472), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n471), .A2(new_n473), .A3(new_n478), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT36), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n397), .A2(KEYINPUT74), .ZN(new_n488));
  INV_X1    g287(.A(new_n393), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT74), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n388), .A2(new_n400), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n388), .A2(KEYINPUT75), .A3(new_n400), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n490), .A2(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n277), .B(new_n278), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n436), .B1(KEYINPUT81), .B2(new_n434), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n444), .B1(new_n499), .B2(new_n439), .ZN(new_n500));
  INV_X1    g299(.A(new_n448), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n450), .A2(new_n487), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n484), .B(new_n485), .C1(new_n500), .C2(new_n501), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n498), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n403), .A2(new_n281), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n479), .A2(new_n480), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT35), .A4(new_n449), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(KEYINPUT84), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n513), .B2(KEYINPUT84), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n514), .A2(new_n517), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n519), .A2(KEYINPUT15), .B1(new_n516), .B2(new_n512), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n532), .B(new_n533), .C1(G1gat), .C2(new_n530), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(G8gat), .Z(new_n535));
  NOR2_X1   g334(.A1(new_n521), .A2(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT17), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n529), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n527), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(KEYINPUT86), .A2(KEYINPUT18), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT88), .B1(new_n539), .B2(new_n527), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n540), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n542), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G197gat), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT11), .B(G169gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT12), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n545), .A2(new_n559), .A3(new_n546), .A4(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n511), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT91), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G155gat), .ZN(new_n565));
  XOR2_X1   g364(.A(G183gat), .B(G211gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n575), .A2(KEYINPUT90), .B1(new_n574), .B2(new_n569), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n575), .A2(KEYINPUT90), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n234), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n234), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n539), .B1(new_n578), .B2(KEYINPUT21), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n581), .A2(new_n234), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n582), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n568), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n585), .B1(new_n583), .B2(new_n584), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n587), .A3(new_n582), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n567), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT41), .ZN(new_n605));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n536), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT94), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n529), .A2(new_n537), .A3(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n605), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT92), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT93), .ZN(new_n615));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n612), .A2(new_n617), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n594), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n578), .B(new_n603), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n455), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT95), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n626), .A2(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n625), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT96), .B(new_n624), .C1(new_n630), .C2(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n562), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n281), .A2(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n281), .A2(KEYINPUT97), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(G1gat), .Z(G1324gat));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n641), .A2(new_n496), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G8gat), .B1(new_n641), .B2(new_n496), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(KEYINPUT98), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n651), .A2(new_n652), .B1(new_n649), .B2(new_n656), .ZN(G1325gat));
  OAI21_X1  g456(.A(G15gat), .B1(new_n641), .B2(new_n487), .ZN(new_n658));
  INV_X1    g457(.A(new_n509), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n641), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT99), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n641), .A2(new_n449), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  AND2_X1   g464(.A1(new_n590), .A2(new_n593), .ZN(new_n666));
  INV_X1    g465(.A(new_n620), .ZN(new_n667));
  INV_X1    g466(.A(new_n638), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n562), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(G29gat), .A3(new_n645), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT100), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n511), .A2(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n504), .A2(new_n676), .A3(new_n507), .A4(new_n510), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n674), .A2(new_n675), .A3(new_n620), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n679), .B(new_n675), .C1(new_n511), .C2(new_n620), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n450), .A2(new_n487), .A3(new_n503), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n507), .A2(new_n510), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n620), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT102), .B1(new_n683), .B2(KEYINPUT44), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n678), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n666), .B(KEYINPUT101), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n561), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n668), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(new_n644), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n673), .B1(new_n522), .B2(new_n691), .ZN(G1328gat));
  NOR3_X1   g491(.A1(new_n670), .A2(G36gat), .A3(new_n496), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT46), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n690), .A2(new_n403), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n523), .ZN(G1329gat));
  INV_X1    g495(.A(new_n487), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n670), .A2(G43gat), .A3(new_n659), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT47), .B1(new_n700), .B2(KEYINPUT104), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n685), .A2(new_n502), .A3(new_n689), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G50gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n449), .A2(G50gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n562), .A2(new_n669), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(KEYINPUT48), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n707), .B(KEYINPUT106), .Z(new_n709));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n704), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n712));
  AOI211_X1 g511(.A(KEYINPUT107), .B(KEYINPUT48), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n705), .A2(new_n710), .ZN(new_n715));
  INV_X1    g514(.A(new_n709), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n708), .B1(new_n713), .B2(new_n719), .ZN(G1331gat));
  AND2_X1   g519(.A1(new_n674), .A2(new_n677), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n594), .A2(new_n620), .A3(new_n638), .A4(new_n561), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n644), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n496), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n723), .B2(new_n487), .ZN(new_n732));
  INV_X1    g531(.A(G71gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n509), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n723), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n735), .B(new_n736), .Z(G1334gat));
  NAND2_X1  g536(.A1(new_n724), .A2(new_n502), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  INV_X1    g538(.A(new_n683), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n666), .A2(new_n561), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n668), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(G85gat), .A3(new_n645), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n666), .A2(new_n561), .A3(new_n638), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n685), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n598), .B1(new_n750), .B2(new_n644), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT109), .ZN(G1336gat));
  NOR3_X1   g552(.A1(new_n747), .A2(G92gat), .A3(new_n496), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n599), .B1(new_n750), .B2(new_n403), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT52), .Z(G1337gat));
  NAND2_X1  g556(.A1(new_n750), .A2(new_n697), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G99gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n638), .A2(G99gat), .A3(new_n659), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n746), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1338gat));
  NAND2_X1  g561(.A1(new_n750), .A2(new_n502), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT53), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n449), .A2(G106gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n747), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n763), .B2(G106gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n766), .B(new_n769), .ZN(G1339gat));
  NOR2_X1   g569(.A1(new_n548), .A2(new_n550), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n541), .A2(new_n542), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n556), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n560), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n668), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n624), .B1(new_n633), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n631), .A2(new_n632), .ZN(new_n778));
  INV_X1    g577(.A(new_n628), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT54), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n778), .A2(new_n779), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n634), .A2(new_n624), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT55), .B(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n785), .A2(new_n561), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n620), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n787), .A2(new_n786), .ZN(new_n790));
  AND4_X1   g589(.A1(new_n620), .A2(new_n790), .A3(new_n774), .A4(new_n785), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n686), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n666), .A2(new_n667), .A3(new_n688), .A4(new_n638), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n621), .A2(new_n795), .A3(new_n688), .A4(new_n638), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n645), .A2(new_n403), .A3(new_n659), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n798), .A2(new_n449), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n688), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n506), .A2(new_n403), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n644), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT113), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n561), .A2(new_n241), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(G1340gat));
  OAI21_X1  g606(.A(G120gat), .B1(new_n801), .B2(new_n638), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n668), .A2(new_n245), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1341gat));
  NAND3_X1  g611(.A1(new_n800), .A2(G127gat), .A3(new_n687), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  INV_X1    g615(.A(new_n804), .ZN(new_n817));
  AOI21_X1  g616(.A(G127gat), .B1(new_n817), .B2(new_n666), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(G1342gat));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n232), .A3(new_n620), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n801), .B2(new_n667), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  NOR2_X1   g623(.A1(new_n697), .A2(new_n449), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n403), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n697), .B2(new_n449), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n645), .B(new_n829), .C1(new_n792), .C2(new_n797), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n561), .A2(new_n205), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT118), .Z(new_n832));
  AOI21_X1  g631(.A(KEYINPUT58), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n644), .A2(new_n496), .A3(new_n487), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT116), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n594), .B1(new_n789), .B2(new_n791), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n797), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n502), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n836), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n798), .A2(new_n841), .A3(new_n502), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n561), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT120), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G141gat), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(KEYINPUT120), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n833), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n848), .A2(new_n842), .A3(new_n835), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n205), .B1(new_n849), .B2(new_n561), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n830), .A2(new_n832), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT119), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT58), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n853), .ZN(G1344gat));
  NAND3_X1  g653(.A1(new_n830), .A2(new_n206), .A3(new_n668), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n798), .A2(KEYINPUT57), .A3(new_n502), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT121), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n667), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n790), .A2(KEYINPUT122), .A3(new_n620), .A4(new_n785), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n774), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n775), .A2(new_n788), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n667), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n666), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n793), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n502), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n841), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n798), .A2(new_n870), .A3(KEYINPUT57), .A4(new_n502), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n858), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n668), .A3(new_n835), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n856), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT59), .B(new_n206), .C1(new_n849), .C2(new_n668), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n855), .B1(new_n874), .B2(new_n875), .ZN(G1345gat));
  INV_X1    g675(.A(new_n849), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n220), .B1(new_n877), .B2(new_n686), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n830), .A2(new_n225), .A3(new_n666), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n877), .B2(new_n667), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n830), .A2(new_n211), .A3(new_n620), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n644), .A2(new_n496), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT123), .Z(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n659), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n798), .A3(new_n449), .ZN(new_n887));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n688), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n798), .A2(new_n884), .ZN(new_n889));
  INV_X1    g688(.A(new_n506), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n561), .A2(new_n324), .A3(new_n325), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1348gat));
  OAI21_X1  g692(.A(new_n283), .B1(new_n891), .B2(new_n638), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT124), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n887), .A2(new_n283), .A3(new_n638), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1349gat));
  OAI21_X1  g696(.A(G183gat), .B1(new_n887), .B2(new_n686), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n666), .A2(new_n292), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n900), .B(new_n901), .Z(G1350gat));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n798), .A3(new_n449), .A4(new_n620), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(G190gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n903), .B2(G190gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n620), .A2(new_n293), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n905), .A2(new_n906), .B1(new_n891), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(G1351gat));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n825), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n561), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n885), .A2(new_n697), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n872), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n561), .A2(G197gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n668), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G204gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n911), .A2(G204gat), .A3(new_n638), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT62), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1353gat));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n355), .A3(new_n666), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n872), .A2(new_n666), .A3(new_n914), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n924), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n924), .B2(G211gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1354gat));
  OAI21_X1  g726(.A(new_n340), .B1(new_n911), .B2(new_n667), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT127), .B(new_n340), .C1(new_n911), .C2(new_n667), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n667), .A2(new_n340), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n915), .B2(new_n933), .ZN(G1355gat));
endmodule


