//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT10), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT65), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n196), .B2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n193), .A3(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n193), .A2(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n196), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n209), .A3(new_n210), .A4(G128), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n192), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT80), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT81), .B1(new_n215), .B2(G104), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n215), .A3(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n213), .A3(G107), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n216), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G101), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT83), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(KEYINPUT79), .A3(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n213), .A2(G107), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n228), .A2(new_n215), .A3(KEYINPUT79), .A4(G104), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n222), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n222), .B2(new_n230), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n212), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT84), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n212), .B(new_n235), .C1(new_n231), .C2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n243), .A3(new_n246), .A4(new_n241), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n247), .A2(new_n248), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n211), .B1(new_n206), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n222), .A2(new_n230), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT82), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n222), .A2(new_n254), .A3(new_n257), .A4(new_n230), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT10), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G101), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n230), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT0), .B(G128), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n198), .B2(new_n202), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n253), .A2(KEYINPUT0), .A3(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n260), .A2(new_n268), .A3(G101), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n262), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n237), .A2(new_n252), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT85), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n237), .A2(KEYINPUT85), .A3(new_n271), .A4(new_n252), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT86), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n237), .A2(new_n271), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n251), .ZN(new_n289));
  INV_X1    g103(.A(new_n284), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n274), .B2(new_n275), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT86), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n231), .A2(new_n232), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n208), .A2(new_n211), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n256), .A2(new_n258), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n251), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n284), .B1(new_n300), .B2(new_n276), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n191), .B1(new_n303), .B2(new_n189), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n190), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n295), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n267), .A2(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G224), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G953), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT7), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n310), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT91), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT2), .B(G113), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G113), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT90), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(new_n320), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n294), .A2(new_n321), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n326), .B1(new_n329), .B2(new_n323), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n321), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n222), .A2(new_n230), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(G110), .B(G122), .Z(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT89), .B(KEYINPUT8), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n316), .B(new_n317), .C1(new_n336), .C2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n294), .A2(new_n321), .A3(new_n332), .ZN(new_n341));
  INV_X1    g155(.A(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n329), .A2(new_n318), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n321), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n262), .A2(new_n344), .A3(new_n269), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n339), .B1(new_n331), .B2(new_n335), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT91), .B1(new_n347), .B2(new_n315), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n345), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n337), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n310), .B(new_n312), .Z(new_n353));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n354), .A3(new_n337), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n356), .A3(new_n189), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n358), .B(KEYINPUT92), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n349), .A2(new_n356), .A3(new_n189), .A4(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G214), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n276), .A2(new_n289), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n290), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n291), .A2(new_n300), .ZN(new_n369));
  AOI21_X1  g183(.A(G902), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n305), .B1(new_n370), .B2(new_n191), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n293), .B2(new_n302), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(new_n191), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT98), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n196), .B2(G128), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n204), .A2(KEYINPUT98), .A3(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT97), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n204), .B2(G143), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n196), .A2(KEYINPUT97), .A3(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n239), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n381), .A3(G134), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n385), .A3(G134), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n386), .A2(new_n382), .ZN(new_n388));
  XNOR2_X1  g202(.A(G116), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT96), .B(G107), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G122), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G116), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n215), .B1(new_n394), .B2(KEYINPUT14), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n389), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n383), .A3(new_n384), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n188), .A2(G217), .A3(new_n277), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n399), .B(KEYINPUT99), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n400), .A3(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n189), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT15), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G478), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n404), .B(new_n189), .C1(KEYINPUT15), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT100), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G237), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n281), .A2(G214), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(new_n196), .ZN(new_n415));
  AOI21_X1  g229(.A(G237), .B1(new_n278), .B2(new_n280), .ZN(new_n416));
  AOI21_X1  g230(.A(G143), .B1(new_n416), .B2(G214), .ZN(new_n417));
  OAI21_X1  g231(.A(G131), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n196), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(G143), .A3(G214), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n246), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G125), .B(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT16), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n307), .A2(G140), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(G146), .C1(KEYINPUT16), .C2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(KEYINPUT16), .B2(new_n426), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n193), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n246), .B1(new_n420), .B2(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n423), .A2(new_n427), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n424), .B(new_n193), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n420), .B(new_n421), .C1(new_n434), .C2(new_n246), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n433), .B(new_n435), .C1(new_n418), .C2(new_n434), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n213), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n432), .A2(new_n436), .A3(new_n439), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n189), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G475), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT93), .B(KEYINPUT20), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT94), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n415), .A2(new_n417), .A3(G131), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n430), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n418), .A2(KEYINPUT94), .A3(new_n422), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n424), .B(KEYINPUT19), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n193), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n427), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n436), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n440), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n442), .ZN(new_n457));
  NOR2_X1   g271(.A1(G475), .A2(G902), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n447), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n460), .A2(KEYINPUT95), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT20), .B1(new_n460), .B2(KEYINPUT95), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n439), .B1(new_n454), .B2(new_n436), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n432), .A2(new_n436), .A3(new_n439), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n445), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G952), .ZN(new_n469));
  AOI211_X1 g283(.A(G953), .B(new_n469), .C1(G234), .C2(G237), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n189), .B(new_n281), .C1(G234), .C2(G237), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT101), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n412), .A2(new_n468), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n306), .A2(new_n366), .A3(new_n373), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n429), .A2(new_n427), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n324), .B2(G128), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n324), .A2(G128), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G110), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT75), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n204), .A2(G119), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT24), .B(G110), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n479), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT76), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n491), .B(new_n492), .C1(G110), .C2(new_n484), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(new_n427), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n491), .B1(new_n484), .B2(G110), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n495), .A2(KEYINPUT76), .B1(new_n193), .B2(new_n424), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT77), .B1(new_n494), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT22), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(G137), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n502), .B(new_n242), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n505), .B(new_n490), .C1(new_n497), .C2(new_n498), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n189), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT25), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n507), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G217), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(G234), .B2(new_n189), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n504), .A2(new_n506), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT66), .B1(new_n264), .B2(new_n266), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT66), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n194), .A2(new_n197), .B1(new_n199), .B2(new_n201), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n518), .B(new_n265), .C1(new_n519), .C2(new_n263), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n251), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n247), .B(new_n248), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n242), .A2(G134), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n246), .B1(new_n241), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n295), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n251), .A2(new_n267), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n526), .A3(KEYINPUT30), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(KEYINPUT68), .A3(new_n528), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n344), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n344), .B(KEYINPUT69), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n536), .A2(new_n532), .A3(new_n526), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n416), .A2(G210), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT26), .B(G101), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n535), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT31), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n535), .A2(new_n546), .A3(new_n538), .A4(new_n543), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n295), .A2(new_n522), .A3(new_n525), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n265), .B1(new_n519), .B2(new_n263), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n522), .B2(new_n245), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n532), .A2(new_n526), .A3(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n536), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n557));
  AOI22_X1  g371(.A1(new_n521), .A2(new_n526), .B1(new_n343), .B2(new_n321), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n537), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n543), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT74), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n563), .B(new_n543), .C1(new_n556), .C2(new_n559), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n545), .B(new_n547), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G472), .A2(G902), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n565), .A2(KEYINPUT32), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT32), .B1(new_n565), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n560), .A2(new_n561), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n543), .B1(new_n535), .B2(new_n538), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT29), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n536), .B1(new_n532), .B2(new_n526), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT28), .B1(new_n537), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n556), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n543), .A2(KEYINPUT29), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n189), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G472), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n516), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n478), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n226), .ZN(G3));
  NAND2_X1  g396(.A1(new_n565), .A2(new_n566), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G472), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n565), .B2(new_n189), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n306), .A2(new_n373), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n516), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n361), .A2(new_n364), .A3(new_n362), .A4(new_n476), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  INV_X1    g405(.A(new_n403), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n400), .B1(new_n392), .B2(new_n397), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n402), .A2(KEYINPUT33), .A3(new_n403), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n594), .A2(new_n595), .A3(G478), .A4(new_n189), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n405), .A2(new_n408), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n600), .B2(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n467), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n590), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n588), .A2(new_n589), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT103), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n604), .B(new_n606), .ZN(G6));
  INV_X1    g421(.A(new_n590), .ZN(new_n608));
  INV_X1    g422(.A(new_n459), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n457), .A2(new_n458), .A3(new_n447), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(G475), .B2(new_n444), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n608), .A2(new_n411), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n588), .A2(new_n589), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G107), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  INV_X1    g429(.A(new_n587), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n617), .A2(new_n499), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n499), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n618), .A2(new_n514), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n510), .B2(new_n512), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n478), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT37), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G110), .ZN(G12));
  AOI21_X1  g440(.A(KEYINPUT86), .B1(new_n276), .B2(new_n284), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n286), .B(new_n290), .C1(new_n274), .C2(new_n275), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n301), .B1(new_n629), .B2(new_n289), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n305), .B(G469), .C1(new_n630), .C2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n190), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n633));
  OR3_X1    g447(.A1(new_n473), .A2(new_n633), .A3(G900), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n473), .B2(G900), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n471), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n611), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n373), .A2(new_n631), .A3(new_n632), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n412), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT32), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n583), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n565), .A2(KEYINPUT32), .A3(new_n566), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n578), .ZN(new_n643));
  INV_X1    g457(.A(new_n621), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n643), .A2(new_n366), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  AND3_X1   g461(.A1(new_n373), .A2(new_n631), .A3(new_n632), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n636), .B(KEYINPUT39), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n648), .A2(KEYINPUT105), .A3(new_n650), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n363), .B(KEYINPUT38), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n644), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n537), .A2(new_n573), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n661), .B2(new_n561), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n535), .A2(new_n538), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n664), .B2(new_n561), .ZN(new_n665));
  AOI211_X1 g479(.A(new_n568), .B(new_n567), .C1(G472), .C2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n365), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n412), .A2(new_n468), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n656), .A2(new_n658), .A3(new_n660), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  NAND3_X1  g485(.A1(new_n601), .A2(new_n467), .A3(new_n636), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n643), .A2(new_n644), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n648), .A2(new_n674), .A3(KEYINPUT106), .A4(new_n366), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n373), .A2(new_n366), .A3(new_n631), .A4(new_n632), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n643), .A2(new_n644), .A3(new_n673), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  AOI22_X1  g495(.A1(new_n367), .A2(new_n290), .B1(new_n291), .B2(new_n300), .ZN(new_n682));
  OAI21_X1  g496(.A(G469), .B1(new_n682), .B2(G902), .ZN(new_n683));
  INV_X1    g497(.A(new_n369), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n284), .B1(new_n276), .B2(new_n289), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n191), .B(new_n189), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n683), .A2(new_n686), .A3(new_n687), .A4(new_n632), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n686), .A3(new_n632), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n579), .A2(new_n603), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT108), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT41), .B(G113), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n579), .A2(new_n612), .A3(new_n688), .A4(new_n690), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AND3_X1   g510(.A1(new_n690), .A2(new_n366), .A3(new_n688), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n621), .B1(new_n569), .B2(new_n578), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n477), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  NOR3_X1   g514(.A1(new_n590), .A2(new_n412), .A3(new_n468), .ZN(new_n701));
  INV_X1    g515(.A(new_n566), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n575), .A2(new_n561), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n547), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n704), .B2(new_n545), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n586), .A2(new_n516), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n701), .A2(new_n690), .A3(new_n688), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  NOR4_X1   g522(.A1(new_n586), .A2(new_n672), .A3(new_n705), .A4(new_n621), .ZN(new_n709));
  AND4_X1   g523(.A1(new_n366), .A2(new_n709), .A3(new_n690), .A4(new_n688), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n307), .ZN(G27));
  AOI21_X1  g525(.A(new_n365), .B1(new_n361), .B2(new_n362), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n632), .ZN(new_n713));
  INV_X1    g527(.A(new_n686), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n293), .A2(KEYINPUT109), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n629), .A2(new_n716), .A3(new_n289), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n301), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n714), .B1(new_n718), .B2(G469), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n191), .A2(new_n189), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n713), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n579), .A3(new_n673), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n716), .B1(new_n629), .B2(new_n289), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n716), .A2(new_n287), .A3(new_n289), .A4(new_n292), .ZN(new_n727));
  OAI211_X1 g541(.A(G469), .B(new_n302), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n686), .A3(new_n721), .ZN(new_n729));
  INV_X1    g543(.A(new_n713), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n579), .A3(new_n673), .A4(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n725), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT111), .B(G131), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G33));
  AND2_X1   g551(.A1(new_n637), .A2(new_n411), .ZN(new_n738));
  AND4_X1   g552(.A1(new_n579), .A2(new_n729), .A3(new_n730), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n239), .ZN(G36));
  NAND2_X1  g554(.A1(new_n718), .A2(KEYINPUT45), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n630), .A2(KEYINPUT45), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(G469), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n721), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT46), .B1(new_n743), .B2(new_n721), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n745), .A3(new_n714), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n190), .A3(new_n649), .ZN(new_n747));
  INV_X1    g561(.A(new_n712), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n468), .A2(new_n601), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT43), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n587), .A3(new_n621), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n748), .B1(new_n751), .B2(KEYINPUT44), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(KEYINPUT44), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n747), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  OAI21_X1  g569(.A(KEYINPUT47), .B1(new_n746), .B2(new_n190), .ZN(new_n756));
  INV_X1    g570(.A(new_n745), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n721), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n686), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n632), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n643), .A2(new_n589), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n748), .A2(new_n672), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n756), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  NAND2_X1  g579(.A1(new_n683), .A2(new_n686), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n632), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n756), .B2(new_n761), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n750), .A2(new_n471), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n706), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n768), .A2(new_n748), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n690), .A2(new_n688), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n748), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n589), .A3(new_n666), .A4(new_n470), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n601), .A2(new_n467), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n774), .A2(new_n769), .ZN(new_n781));
  OR4_X1    g595(.A1(new_n586), .A2(new_n781), .A3(new_n621), .A4(new_n705), .ZN(new_n782));
  INV_X1    g596(.A(new_n657), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n773), .A2(KEYINPUT115), .A3(new_n364), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT115), .B1(new_n773), .B2(new_n364), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(KEYINPUT50), .A3(new_n770), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT50), .B1(new_n786), .B2(new_n770), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n780), .B(new_n782), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n772), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n756), .A2(new_n761), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n712), .B(new_n770), .C1(new_n791), .C2(new_n767), .ZN(new_n792));
  INV_X1    g606(.A(new_n789), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n410), .B(KEYINPUT112), .Z(new_n797));
  NOR2_X1   g611(.A1(new_n748), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n643), .A3(new_n644), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n638), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n739), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n722), .A2(new_n802), .A3(new_n709), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n729), .A2(new_n709), .A3(new_n730), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT113), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n735), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n710), .B1(new_n639), .B2(new_n645), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n621), .A2(new_n636), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n809), .A2(new_n363), .A3(new_n190), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n667), .A2(new_n668), .A3(new_n729), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n680), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n699), .A2(new_n691), .A3(new_n695), .A4(new_n707), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n306), .A2(new_n373), .A3(new_n587), .ZN(new_n816));
  INV_X1    g630(.A(new_n602), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n468), .B2(new_n797), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n816), .A2(new_n516), .A3(new_n590), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n478), .B1(new_n580), .B2(new_n623), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n815), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n680), .A2(new_n808), .A3(new_n811), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n807), .A2(new_n814), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n735), .A2(new_n801), .A3(new_n806), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n695), .A2(new_n691), .A3(new_n707), .ZN(new_n828));
  INV_X1    g642(.A(new_n818), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n588), .A2(new_n589), .A3(new_n608), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n677), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(new_n477), .C1(new_n579), .C2(new_n622), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n699), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n680), .A2(new_n808), .A3(new_n811), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n826), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n807), .A2(new_n821), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n836), .A2(new_n838), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT53), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n834), .A2(new_n835), .A3(new_n814), .A4(new_n824), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n781), .A2(new_n580), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT48), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n777), .A2(new_n817), .A3(new_n778), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(G952), .A3(new_n277), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n697), .B2(new_n770), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n842), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT117), .B1(new_n796), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n469), .A2(new_n277), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n790), .A2(new_n795), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n845), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT54), .B1(new_n826), .B2(new_n839), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n859), .A3(new_n860), .A4(new_n852), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n854), .A2(new_n855), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n783), .B1(new_n766), .B2(KEYINPUT49), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n749), .A2(new_n516), .A3(new_n365), .A4(new_n190), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n766), .A2(KEYINPUT49), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n666), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n862), .A2(new_n866), .ZN(G75));
  NAND2_X1  g681(.A1(new_n352), .A2(new_n355), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n353), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT55), .Z(new_n870));
  NAND3_X1  g684(.A1(new_n826), .A2(G902), .A3(new_n839), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n360), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n872), .B2(KEYINPUT56), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n281), .A2(G952), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT120), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n826), .A2(new_n839), .A3(new_n880), .A4(G902), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n882), .B2(new_n359), .ZN(new_n883));
  AOI211_X1 g697(.A(KEYINPUT119), .B(new_n360), .C1(new_n879), .C2(new_n881), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(G51));
  XNOR2_X1  g701(.A(new_n720), .B(KEYINPUT57), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n826), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n858), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n685), .B2(new_n684), .ZN(new_n891));
  INV_X1    g705(.A(new_n743), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n874), .B1(new_n891), .B2(new_n893), .ZN(G54));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n879), .B2(new_n881), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n896), .A2(G475), .A3(new_n457), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n457), .B1(new_n896), .B2(G475), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n874), .ZN(G60));
  NAND2_X1  g713(.A1(new_n594), .A2(new_n595), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n901), .B(new_n904), .C1(new_n889), .C2(new_n858), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n842), .B2(new_n847), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n907), .B2(new_n901), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n909), .B(new_n900), .C1(new_n859), .C2(new_n903), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n875), .B(new_n906), .C1(new_n908), .C2(new_n910), .ZN(G63));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n826), .A2(new_n839), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n504), .A2(new_n506), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n875), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n618), .A2(new_n619), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n826), .A2(new_n839), .A3(new_n918), .A4(new_n914), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(KEYINPUT61), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT61), .B1(new_n917), .B2(new_n919), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n926), .B(KEYINPUT61), .C1(new_n917), .C2(new_n919), .ZN(new_n927));
  OAI22_X1  g741(.A1(new_n922), .A2(new_n923), .B1(new_n925), .B2(new_n927), .ZN(G66));
  INV_X1    g742(.A(new_n281), .ZN(new_n929));
  INV_X1    g743(.A(new_n475), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n930), .B2(new_n311), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n821), .A2(new_n929), .B1(KEYINPUT124), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(KEYINPUT124), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n868), .B1(G898), .B2(new_n281), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(G69));
  AOI21_X1  g749(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n452), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(G900), .B2(new_n929), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n366), .A2(new_n668), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n747), .A2(new_n942), .A3(new_n579), .A4(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n759), .A2(new_n579), .A3(new_n632), .A4(new_n650), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT126), .B1(new_n946), .B2(new_n943), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n680), .A2(new_n808), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n735), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n739), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n764), .A2(new_n754), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n941), .B1(new_n953), .B2(new_n281), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n764), .A2(new_n754), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n945), .A2(new_n947), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n958), .A3(new_n951), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n940), .B1(new_n959), .B2(new_n929), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT127), .B1(new_n960), .B2(KEYINPUT125), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n936), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n670), .A2(new_n949), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n655), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(new_n579), .A3(new_n712), .A4(new_n829), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n965), .A2(new_n957), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n938), .B1(new_n968), .B2(new_n929), .ZN(new_n969));
  INV_X1    g783(.A(new_n936), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n969), .A2(KEYINPUT125), .A3(new_n970), .A4(new_n960), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n962), .A2(new_n971), .ZN(G72));
  NAND4_X1  g786(.A1(new_n965), .A2(new_n821), .A3(new_n957), .A4(new_n967), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n664), .A2(new_n561), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n874), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n571), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n544), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n845), .A2(new_n846), .A3(new_n975), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n975), .B1(new_n959), .B2(new_n833), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n664), .A3(new_n561), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(G57));
endmodule


