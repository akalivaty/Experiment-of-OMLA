//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n214), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n250), .B(new_n251), .C1(new_n252), .C2(new_n248), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n208), .A2(G274), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT66), .B(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n261), .B1(G226), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G200), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n267));
  INV_X1    g0067(.A(G150), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n267), .B1(new_n268), .B2(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n215), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n209), .A2(G1), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n201), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n281), .A2(new_n283), .B1(new_n201), .B2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT9), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n257), .A2(G190), .A3(new_n264), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n278), .A2(KEYINPUT9), .A3(new_n284), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n266), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT10), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(KEYINPUT10), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n265), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n257), .A2(new_n296), .A3(new_n264), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n285), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT66), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G45), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n308), .A3(new_n260), .ZN(new_n309));
  INV_X1    g0109(.A(new_n258), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n255), .A2(G238), .A3(new_n262), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n249), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n232), .A2(G1698), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n255), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT13), .B1(new_n313), .B2(new_n321), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G190), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT75), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(KEYINPUT74), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT74), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(KEYINPUT13), .C1(new_n313), .C2(new_n321), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT73), .B1(new_n322), .B2(new_n323), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  NOR4_X1   g0132(.A1(new_n313), .A2(new_n321), .A3(new_n332), .A4(KEYINPUT13), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n273), .A2(new_n252), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n270), .A2(new_n201), .B1(new_n209), .B2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n277), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n339), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n280), .A2(new_n220), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT12), .ZN(new_n343));
  INV_X1    g0143(.A(new_n282), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n281), .A2(G68), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(new_n341), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n327), .A2(new_n335), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n277), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n274), .A2(new_n270), .B1(new_n209), .B2(new_n252), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT70), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT70), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n356), .A3(new_n272), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n350), .B1(new_n357), .B2(KEYINPUT71), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT71), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n353), .A2(new_n356), .A3(new_n359), .A4(new_n272), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n349), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n281), .A2(G77), .A3(new_n344), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G77), .B2(new_n279), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n263), .A2(G244), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n311), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G238), .A2(G1698), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n232), .B2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n248), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G107), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G107), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n369), .B1(new_n248), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n255), .B1(new_n375), .B2(KEYINPUT69), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT69), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n369), .B(new_n377), .C1(new_n248), .C2(new_n374), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n366), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G190), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n364), .B(new_n380), .C1(new_n381), .C2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n348), .A2(new_n382), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n361), .A2(new_n363), .B1(new_n379), .B2(G169), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(KEYINPUT72), .B1(new_n296), .B2(new_n379), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT72), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n386), .B1(new_n379), .B2(G169), .C1(new_n361), .C2(new_n363), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n304), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n314), .A2(G1698), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G223), .B2(G1698), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n317), .A2(new_n318), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n271), .B2(new_n222), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n261), .B1(new_n393), .B2(new_n256), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n255), .A2(G232), .A3(new_n262), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT76), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n255), .A2(new_n262), .A3(new_n397), .A4(G232), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n381), .ZN(new_n401));
  INV_X1    g0201(.A(G190), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n392), .B2(new_n209), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n317), .A2(new_n318), .A3(new_n407), .A4(G20), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n202), .A2(new_n220), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n269), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n405), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(KEYINPUT3), .A2(G33), .ZN(new_n417));
  NAND2_X1  g0217(.A1(KEYINPUT3), .A2(G33), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n209), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n407), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n417), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n418), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n220), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n277), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n281), .ZN(new_n425));
  INV_X1    g0225(.A(new_n274), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n344), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n425), .A2(new_n427), .B1(new_n426), .B2(new_n279), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n404), .A2(new_n424), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT16), .B1(new_n422), .B2(new_n414), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n409), .A2(new_n405), .A3(new_n415), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n428), .B1(new_n435), .B2(new_n277), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n400), .A2(new_n294), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G179), .B2(new_n400), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT18), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n394), .A2(new_n296), .A3(new_n399), .ZN(new_n440));
  AOI21_X1  g0240(.A(G169), .B1(new_n394), .B2(new_n399), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n349), .B1(new_n433), .B2(new_n434), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n428), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n404), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n432), .A2(new_n439), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n324), .A2(G179), .A3(new_n325), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n334), .A2(KEYINPUT14), .A3(G169), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT14), .B1(new_n334), .B2(G169), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n447), .B1(new_n452), .B2(new_n346), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n389), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n209), .B(G87), .C1(new_n317), .C2(new_n318), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT22), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT22), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n248), .A2(new_n457), .A3(new_n209), .A4(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n370), .A2(G20), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(KEYINPUT23), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n371), .A2(new_n373), .A3(G20), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(KEYINPUT23), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT24), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n467), .A3(new_n464), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n349), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G13), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n461), .A2(G1), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n208), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n279), .A2(new_n474), .A3(new_n215), .A4(new_n276), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n370), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT83), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n468), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n467), .B1(new_n459), .B2(new_n464), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n277), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n477), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n485));
  OAI211_X1 g0285(.A(G250), .B(new_n249), .C1(new_n317), .C2(new_n318), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT84), .A2(G294), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT84), .A2(G294), .ZN(new_n488));
  OAI21_X1  g0288(.A(G33), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n256), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n208), .A2(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G274), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT5), .B(G41), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n305), .A2(G1), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n498), .A2(new_n499), .B1(new_n216), .B2(new_n254), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G264), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G169), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n490), .A2(new_n256), .B1(new_n500), .B2(G264), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G179), .A3(new_n497), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n479), .A2(new_n484), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n381), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(G190), .B2(new_n502), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n482), .A3(new_n477), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  MUX2_X1   g0311(.A(new_n279), .B(new_n475), .S(G116), .Z(new_n512));
  INV_X1    g0312(.A(G116), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G20), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n277), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n516));
  AOI21_X1  g0316(.A(G20), .B1(G33), .B2(G283), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n271), .A2(G97), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT80), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT80), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n515), .B(new_n516), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT81), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n277), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n517), .A2(new_n518), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT80), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n528), .B2(new_n519), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n512), .B(new_n522), .C1(new_n524), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(new_n249), .C1(new_n317), .C2(new_n318), .ZN(new_n533));
  XNOR2_X1  g0333(.A(KEYINPUT79), .B(G303), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n248), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n256), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n500), .A2(G270), .B1(G274), .B2(new_n496), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT21), .A3(G169), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(G179), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n531), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n536), .A2(new_n537), .A3(G190), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n381), .B1(new_n536), .B2(new_n537), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n542), .A2(new_n543), .A3(new_n530), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n294), .B1(new_n536), .B2(new_n537), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT21), .B1(new_n545), .B2(new_n530), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n541), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n279), .B1(new_n353), .B2(new_n356), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n475), .A2(new_n222), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G87), .A2(G97), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n371), .A2(new_n373), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n209), .B1(new_n320), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n209), .B(G68), .C1(new_n317), .C2(new_n318), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n552), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(KEYINPUT78), .A3(new_n553), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n548), .B(new_n549), .C1(new_n562), .C2(new_n277), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n221), .A2(new_n249), .ZN(new_n564));
  INV_X1    g0364(.A(G244), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G1698), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n566), .C1(new_n317), .C2(new_n318), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n567), .A2(KEYINPUT77), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT77), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(new_n255), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n499), .A2(new_n223), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n255), .B1(G45), .B2(new_n310), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n567), .A2(new_n568), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT77), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n255), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n567), .A2(KEYINPUT77), .A3(new_n568), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n563), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n294), .B1(new_n571), .B2(new_n574), .ZN(new_n583));
  INV_X1    g0383(.A(new_n548), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n353), .A2(new_n356), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n585), .A2(new_n475), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n551), .A2(KEYINPUT78), .A3(new_n553), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT78), .B1(new_n551), .B2(new_n553), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n557), .A2(new_n559), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n584), .B(new_n586), .C1(new_n590), .C2(new_n349), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n576), .A2(new_n577), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n256), .A3(new_n579), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n296), .A3(new_n573), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n583), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n582), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G244), .B(new_n249), .C1(new_n317), .C2(new_n318), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G283), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n271), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G250), .A2(G1698), .ZN(new_n602));
  NAND2_X1  g0402(.A1(KEYINPUT4), .A2(G244), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(G1698), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n248), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n255), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n495), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n499), .B1(new_n607), .B2(new_n493), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(G257), .A3(new_n255), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n497), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n296), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n294), .B1(new_n606), .B2(new_n610), .ZN(new_n613));
  INV_X1    g0413(.A(new_n374), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n406), .B2(new_n408), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  AND2_X1   g0416(.A1(G97), .A2(G107), .ZN(new_n617));
  NOR2_X1   g0417(.A1(G97), .A2(G107), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n370), .A2(KEYINPUT6), .A3(G97), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n349), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G97), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n280), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n475), .B2(new_n624), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n612), .B(new_n613), .C1(new_n623), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n615), .A2(new_n622), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n628), .B2(new_n277), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n606), .A2(new_n610), .A3(G190), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n599), .A2(new_n605), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n256), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n497), .A2(new_n609), .ZN(new_n633));
  AOI21_X1  g0433(.A(G200), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n547), .A2(new_n596), .A3(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n454), .A2(new_n511), .A3(new_n637), .ZN(G372));
  AND2_X1   g0438(.A1(new_n439), .A2(new_n445), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n448), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n331), .A2(new_n333), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n328), .A2(new_n330), .ZN(new_n643));
  OAI21_X1  g0443(.A(G169), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n641), .B1(new_n646), .B2(new_n449), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n327), .A2(new_n335), .A3(new_n347), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n385), .A2(new_n387), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n347), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n404), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT17), .B1(new_n436), .B2(new_n404), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n640), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n293), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n303), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n454), .ZN(new_n658));
  AOI21_X1  g0458(.A(G169), .B1(new_n632), .B2(new_n633), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n606), .A2(new_n610), .A3(G179), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n629), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n582), .A3(new_n595), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n661), .A2(new_n582), .A3(KEYINPUT26), .A4(new_n595), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n506), .B1(new_n469), .B2(new_n478), .ZN(new_n667));
  INV_X1    g0467(.A(new_n546), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT21), .ZN(new_n669));
  AOI211_X1 g0469(.A(new_n669), .B(new_n294), .C1(new_n536), .C2(new_n537), .ZN(new_n670));
  INV_X1    g0470(.A(new_n540), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n530), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n596), .A3(new_n510), .A4(new_n636), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n666), .A2(new_n674), .A3(new_n595), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n658), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n657), .A2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n530), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n547), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n541), .A2(new_n546), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n479), .A2(new_n484), .A3(new_n683), .ZN(new_n690));
  INV_X1    g0490(.A(new_n683), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n511), .A2(new_n690), .B1(new_n507), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n667), .A2(new_n683), .ZN(new_n694));
  INV_X1    g0494(.A(new_n511), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n686), .A2(new_n683), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(G399));
  NOR2_X1   g0498(.A1(new_n551), .A2(G116), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT85), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n212), .A2(new_n260), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n218), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n611), .A2(new_n504), .A3(new_n593), .A4(new_n573), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n540), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n504), .A2(new_n632), .A3(new_n633), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n671), .A3(KEYINPUT30), .A4(new_n580), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n611), .A2(G179), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n593), .A2(new_n573), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n502), .A3(new_n538), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n708), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n683), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n582), .A2(new_n627), .A3(new_n595), .A4(new_n635), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n695), .A2(new_n722), .A3(new_n547), .A4(new_n691), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n705), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n595), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n664), .B2(new_n665), .ZN(new_n726));
  INV_X1    g0526(.A(new_n510), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n507), .A2(new_n686), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT86), .B1(new_n731), .B2(new_n691), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT86), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n733), .B(new_n683), .C1(new_n726), .C2(new_n730), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT29), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n683), .B1(new_n726), .B2(new_n674), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n724), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n704), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n470), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n208), .B1(new_n740), .B2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n701), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n212), .A2(new_n248), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n744), .A2(new_n206), .B1(G116), .B2(new_n212), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n243), .A2(new_n305), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n212), .A2(new_n392), .ZN(new_n747));
  INV_X1    g0547(.A(new_n218), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(new_n259), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n215), .B1(G20), .B2(new_n294), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n743), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n402), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n209), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n487), .A2(new_n488), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n392), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G20), .A2(G179), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT88), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n402), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(new_n402), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n209), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT89), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT89), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n761), .B(new_n772), .C1(G303), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n402), .A3(G200), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n773), .A2(new_n402), .A3(new_n381), .ZN(new_n781));
  INV_X1    g0581(.A(G329), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n780), .A2(new_n600), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n763), .A2(G190), .A3(new_n381), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(KEYINPUT91), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(KEYINPUT91), .B2(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT90), .Z(new_n791));
  OAI211_X1 g0591(.A(new_n779), .B(new_n788), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n778), .A2(G87), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n201), .B2(new_n790), .C1(new_n252), .C2(new_n770), .ZN(new_n794));
  INV_X1    g0594(.A(new_n781), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n780), .A2(new_n370), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n248), .B1(new_n759), .B2(new_n624), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n786), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G58), .A2(new_n801), .B1(new_n765), .B2(G68), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n792), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n757), .B1(new_n804), .B2(new_n754), .ZN(new_n805));
  INV_X1    g0605(.A(new_n753), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n687), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n687), .A2(G330), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT87), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n688), .A2(new_n742), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(G396));
  OAI21_X1  g0611(.A(new_n683), .B1(new_n361), .B2(new_n363), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n385), .A2(new_n387), .B1(new_n382), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n376), .A2(new_n378), .ZN(new_n814));
  INV_X1    g0614(.A(new_n366), .ZN(new_n815));
  AOI21_X1  g0615(.A(G169), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT72), .B1(new_n364), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n379), .A2(new_n296), .ZN(new_n818));
  AND4_X1   g0618(.A1(new_n387), .A2(new_n817), .A3(new_n812), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n736), .B(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n724), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n743), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  INV_X1    g0624(.A(new_n754), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n752), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n743), .B1(new_n826), .B2(G77), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G159), .A2(new_n769), .B1(new_n801), .B2(G143), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n829), .B2(new_n790), .C1(new_n268), .C2(new_n764), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n392), .B1(new_n795), .B2(G132), .ZN(new_n832));
  INV_X1    g0632(.A(new_n780), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G68), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n834), .C1(new_n202), .C2(new_n759), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G50), .B2(new_n778), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n392), .B1(new_n777), .B2(new_n370), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT93), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n833), .A2(G87), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n840), .B1(new_n624), .B2(new_n759), .C1(new_n771), .C2(new_n781), .ZN(new_n841));
  XOR2_X1   g0641(.A(KEYINPUT92), .B(G283), .Z(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n765), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n769), .A2(G116), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G294), .A2(new_n801), .B1(new_n846), .B2(G303), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n837), .B1(new_n839), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n827), .B1(new_n849), .B2(new_n754), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n752), .B2(new_n820), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n824), .A2(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n621), .A2(KEYINPUT35), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n853), .A2(new_n513), .A3(new_n217), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(KEYINPUT94), .B1(KEYINPUT35), .B2(new_n621), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(KEYINPUT94), .B2(new_n855), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT36), .Z(new_n858));
  OAI211_X1 g0658(.A(new_n748), .B(G77), .C1(new_n202), .C2(new_n220), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n201), .A2(G68), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n208), .B(G13), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  INV_X1    g0663(.A(new_n681), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n444), .B2(new_n428), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n639), .B2(new_n653), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n865), .B2(KEYINPUT96), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n442), .B1(new_n444), .B2(new_n428), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n430), .A4(new_n865), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n681), .B1(new_n424), .B2(new_n429), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT96), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n430), .A3(new_n865), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n863), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n447), .A2(new_n871), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n875), .A4(new_n870), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n675), .A2(new_n820), .A3(new_n691), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n388), .A2(new_n691), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT95), .B1(new_n647), .B2(new_n347), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT95), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n452), .A2(new_n885), .A3(new_n346), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n347), .A2(new_n691), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n648), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n452), .B2(new_n648), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n880), .A2(new_n883), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n639), .A2(new_n864), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n877), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n867), .B1(new_n865), .B2(KEYINPUT98), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n897), .A2(new_n869), .A3(new_n430), .A4(new_n865), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT98), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n871), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n874), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n863), .B1(new_n866), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT39), .B1(new_n903), .B2(new_n879), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n884), .A2(new_n886), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n683), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n895), .A2(KEYINPUT97), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n881), .A2(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n893), .B1(new_n909), .B2(new_n880), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT97), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n454), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n656), .B1(new_n735), .B2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n913), .B(new_n916), .Z(new_n917));
  OR2_X1    g0717(.A1(new_n813), .A2(new_n819), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n720), .B2(new_n723), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n880), .A2(new_n891), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n891), .A2(new_n919), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n903), .B2(new_n879), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n637), .A2(new_n511), .A3(new_n683), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n658), .B1(new_n927), .B2(new_n719), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(G330), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n917), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n208), .B2(new_n740), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n917), .A2(new_n931), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n862), .B1(new_n933), .B2(new_n934), .ZN(G367));
  OAI211_X1 g0735(.A(new_n627), .B(new_n635), .C1(new_n629), .C2(new_n691), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n627), .B2(new_n691), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n695), .A2(new_n696), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n627), .B1(new_n507), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n691), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT99), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n563), .A2(new_n691), .ZN(new_n945));
  MUX2_X1   g0745(.A(new_n596), .B(new_n725), .S(new_n945), .Z(new_n946));
  NOR3_X1   g0746(.A1(new_n944), .A2(KEYINPUT43), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n946), .B(KEYINPUT43), .Z(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n693), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n937), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n701), .B(KEYINPUT41), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n697), .A2(new_n694), .A3(new_n937), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT45), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n937), .B1(new_n697), .B2(new_n694), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT44), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n693), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT100), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n950), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n697), .B1(new_n692), .B2(new_n696), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n689), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n738), .A2(KEYINPUT101), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n738), .A2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT101), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n960), .A2(KEYINPUT100), .A3(new_n950), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n962), .A2(new_n965), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n953), .B1(new_n970), .B2(new_n738), .ZN(new_n971));
  INV_X1    g0771(.A(new_n741), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n952), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n755), .B1(new_n212), .B2(new_n585), .C1(new_n238), .C2(new_n747), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(new_n743), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n392), .B1(new_n795), .B2(G137), .ZN(new_n976));
  INV_X1    g0776(.A(new_n759), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(G68), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n833), .A2(G77), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G150), .A2(new_n801), .B1(new_n765), .B2(G159), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n202), .B2(new_n777), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(G50), .C2(new_n769), .ZN(new_n983));
  INV_X1    g0783(.A(G143), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(new_n791), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT104), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n780), .A2(new_n624), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n248), .B(new_n988), .C1(G317), .C2(new_n795), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT103), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n374), .B2(new_n759), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n989), .A2(KEYINPUT103), .B1(new_n760), .B2(new_n764), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n770), .A2(new_n842), .B1(new_n534), .B2(new_n786), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n791), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT102), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n777), .B2(new_n513), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n995), .A2(G311), .B1(KEYINPUT46), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n994), .B(new_n998), .C1(KEYINPUT46), .C2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n987), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT47), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n754), .B1(new_n1001), .B2(KEYINPUT47), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n975), .B1(new_n806), .B2(new_n946), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n973), .A2(new_n1005), .ZN(G387));
  NAND2_X1  g0806(.A1(new_n426), .A2(new_n201), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n1008), .C1(G68), .C2(G77), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n747), .B1(new_n1009), .B2(new_n700), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n259), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n235), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT105), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(G107), .B2(new_n212), .C1(new_n700), .C2(new_n744), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n742), .B1(new_n1015), .B2(new_n755), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n585), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n977), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT106), .B(G150), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n392), .B1(new_n795), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n624), .C2(new_n780), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G50), .A2(new_n801), .B1(new_n765), .B2(new_n426), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n220), .B2(new_n770), .C1(new_n252), .C2(new_n777), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(G159), .C2(new_n846), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G311), .A2(new_n765), .B1(new_n801), .B2(G317), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n534), .B2(new_n770), .C1(new_n791), .C2(new_n785), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n777), .A2(new_n760), .B1(new_n759), .B2(new_n842), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT49), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT107), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n392), .B1(new_n781), .B2(new_n789), .C1(new_n513), .C2(new_n780), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1032), .B2(KEYINPUT107), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1024), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1016), .B1(new_n692), .B2(new_n806), .C1(new_n1036), .C2(new_n825), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n964), .A2(new_n972), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n966), .A2(new_n260), .A3(new_n212), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n738), .A2(new_n964), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1038), .C1(new_n1039), .C2(new_n1040), .ZN(G393));
  OAI221_X1 g0841(.A(new_n755), .B1(new_n624), .B2(new_n212), .C1(new_n246), .C2(new_n747), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n743), .ZN(new_n1043));
  INV_X1    g0843(.A(G159), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n268), .A2(new_n790), .B1(new_n786), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT51), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n765), .A2(G50), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n977), .A2(G77), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n392), .B1(new_n795), .B2(G143), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1047), .A2(new_n840), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n770), .A2(new_n274), .B1(new_n220), .B2(new_n777), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1046), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT108), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT108), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G311), .A2(new_n801), .B1(new_n846), .B2(G317), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT52), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n248), .B(new_n798), .C1(G322), .C2(new_n795), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n513), .B2(new_n759), .C1(new_n534), .C2(new_n764), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n769), .A2(G294), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n777), .B2(new_n842), .ZN(new_n1060));
  OR3_X1    g0860(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1053), .A2(new_n1054), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1043), .B1(new_n1062), .B2(new_n754), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n806), .B2(new_n937), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n961), .A2(new_n958), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n741), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n701), .B1(new_n1065), .B2(new_n966), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n970), .B2(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT109), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT109), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(G390));
  OAI22_X1  g0871(.A1(new_n909), .A2(new_n907), .B1(new_n896), .B2(new_n904), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n891), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n820), .B1(new_n732), .B2(new_n734), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n882), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n903), .A2(new_n879), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n683), .B2(new_n906), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1072), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n891), .A2(new_n919), .A3(G330), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1072), .B(new_n1079), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n972), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n743), .B1(new_n826), .B2(new_n426), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n778), .A2(new_n1019), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(KEYINPUT53), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1085), .A2(KEYINPUT53), .ZN(new_n1087));
  INV_X1    g0887(.A(G132), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n786), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n392), .B1(new_n795), .B2(G125), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n201), .B2(new_n780), .C1(new_n1044), .C2(new_n759), .ZN(new_n1091));
  OR4_X1    g0891(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n846), .A2(G128), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT54), .B(G143), .Z(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT111), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1093), .B1(new_n829), .B2(new_n764), .C1(new_n770), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n248), .B1(new_n795), .B2(G294), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n793), .A2(new_n834), .A3(new_n1048), .A4(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G97), .A2(new_n769), .B1(new_n846), .B2(G283), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n513), .B2(new_n786), .C1(new_n374), .C2(new_n764), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1092), .A2(new_n1096), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n754), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n905), .B2(new_n752), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n735), .A2(new_n915), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n658), .A2(new_n724), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n657), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT110), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n820), .B1(new_n927), .B2(new_n719), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n889), .B(new_n890), .C1(new_n1110), .C2(new_n705), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1079), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n883), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1079), .A2(new_n1074), .A3(new_n882), .A4(new_n1111), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT110), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n916), .A2(new_n1116), .A3(new_n1107), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1109), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n701), .B1(new_n1105), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(new_n1081), .A3(new_n1082), .A4(new_n1115), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1104), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(new_n1115), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1105), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT115), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n293), .A2(new_n298), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n681), .B1(new_n278), .B2(new_n284), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1128), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n293), .A2(new_n298), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1132), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1130), .B1(new_n293), .B2(new_n298), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1128), .B(new_n299), .C1(new_n291), .C2(new_n292), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1110), .B1(new_n889), .B2(new_n890), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n705), .B1(new_n1139), .B2(new_n924), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n1140), .B2(new_n922), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1133), .A2(new_n1137), .A3(KEYINPUT114), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT114), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1140), .A2(new_n922), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n913), .B(new_n1126), .C1(new_n1141), .C2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n877), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1076), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n907), .B(new_n1147), .C1(new_n1148), .C2(KEYINPUT39), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n910), .B2(new_n911), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n895), .A2(KEYINPUT97), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1145), .A2(new_n1141), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1138), .ZN(new_n1153));
  OAI21_X1  g0953(.A(G330), .B1(new_n925), .B2(new_n923), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT40), .B1(new_n1139), .B2(new_n880), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1140), .A2(new_n922), .A3(new_n1144), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1156), .A2(new_n908), .A3(new_n912), .A4(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(new_n1158), .A3(KEYINPUT115), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1125), .A2(new_n1146), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n701), .B1(new_n1125), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n972), .A3(new_n1146), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n743), .B1(new_n826), .B2(G50), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n248), .A2(G41), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G283), .B2(new_n795), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n978), .C1(new_n202), .C2(new_n780), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G77), .B2(new_n778), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n786), .A2(new_n370), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT112), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n765), .A2(G97), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1017), .A2(new_n769), .B1(new_n846), .B2(G116), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G50), .B1(new_n271), .B2(new_n260), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n1169), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G125), .A2(new_n846), .B1(new_n801), .B2(G128), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n1088), .B2(new_n764), .C1(new_n829), .C2(new_n770), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n777), .A2(new_n1095), .B1(new_n268), .B2(new_n759), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT113), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1044), .C2(new_n780), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1185), .A2(KEYINPUT113), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1180), .B1(new_n1178), .B2(new_n1177), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1167), .B1(new_n1190), .B2(new_n754), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1144), .B2(new_n752), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1166), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1165), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT116), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1124), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n953), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n1118), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1073), .A2(new_n751), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n743), .B1(new_n826), .B2(G68), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n248), .B1(new_n795), .B2(G303), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1018), .A2(new_n979), .A3(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n778), .A2(G97), .B1(G283), .B2(new_n801), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n765), .A2(G116), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n614), .A2(new_n769), .B1(new_n846), .B2(G294), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1095), .A2(new_n764), .B1(new_n1088), .B2(new_n790), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G137), .B2(new_n801), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT117), .Z(new_n1213));
  AOI22_X1  g1013(.A1(new_n977), .A2(G50), .B1(new_n795), .B2(G128), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n777), .B2(new_n1044), .C1(new_n770), .C2(new_n268), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n248), .B1(new_n780), .B2(new_n202), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT118), .Z(new_n1217));
  OR2_X1    g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1210), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT119), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n825), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1204), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1115), .A2(new_n972), .B1(new_n1203), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1202), .A2(new_n1224), .ZN(G381));
  NAND4_X1  g1025(.A1(new_n973), .A2(new_n1005), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1226));
  OR2_X1    g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  OR3_X1    g1027(.A1(G381), .A2(new_n1227), .A3(G384), .ZN(new_n1228));
  OR4_X1    g1028(.A1(G378), .A2(G375), .A3(new_n1226), .A4(new_n1228), .ZN(G407));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1197), .A2(new_n1122), .A3(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT120), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(G407), .A2(new_n1233), .A3(G213), .ZN(G409));
  NAND2_X1  g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1227), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(G387), .A2(G390), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1226), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1238), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G387), .A2(G390), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1238), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1244), .A2(new_n1226), .A3(new_n1245), .A4(new_n1240), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1242), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT121), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1122), .B(new_n1193), .C1(new_n1162), .C2(new_n1164), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1125), .A2(new_n1201), .A3(new_n1146), .A4(new_n1159), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1192), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n972), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1122), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1248), .B1(new_n1249), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1231), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1165), .A2(G378), .A3(new_n1194), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1255), .A3(KEYINPUT121), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n701), .B1(new_n1262), .B2(new_n1200), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1200), .B2(new_n1262), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G384), .B(KEYINPUT122), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1224), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1231), .A2(G2897), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1264), .A2(new_n1224), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1266), .B(new_n1267), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1266), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1270), .B1(new_n1264), .B2(new_n1224), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G2897), .B(new_n1231), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1261), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1257), .A2(new_n1258), .A3(new_n1276), .A4(new_n1260), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1231), .B1(new_n1259), .B2(new_n1255), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1247), .A2(new_n1275), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1242), .A2(KEYINPUT126), .A3(new_n1246), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT126), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1274), .A2(new_n1271), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1243), .B1(new_n1286), .B2(new_n1280), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1277), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1280), .A2(KEYINPUT62), .A3(new_n1276), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI211_X1 g1093(.A(KEYINPUT125), .B(new_n1287), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1282), .B1(new_n1293), .B2(new_n1294), .ZN(G405));
  OAI21_X1  g1095(.A(new_n1259), .B1(new_n1197), .B2(G378), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1276), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  OAI221_X1 g1099(.A(new_n1259), .B1(KEYINPUT127), .B2(new_n1297), .C1(new_n1197), .C2(G378), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1285), .ZN(G402));
endmodule


