//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n188), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT64), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n191), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT66), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G134), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT65), .A3(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT11), .B1(new_n205), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n203), .A3(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n201), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  AND4_X1   g027(.A1(new_n212), .A2(new_n204), .A3(new_n206), .A4(new_n201), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n200), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n217));
  INV_X1    g031(.A(G113), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n219), .A2(new_n220), .B1(KEYINPUT2), .B2(G113), .ZN(new_n221));
  XNOR2_X1  g035(.A(G116), .B(G119), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n196), .A2(G128), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n193), .B(new_n195), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n212), .A2(new_n230), .A3(new_n204), .A4(new_n206), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g046(.A(G134), .B(G137), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n203), .A2(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n205), .A2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT67), .A3(G131), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n229), .A2(new_n231), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n215), .A2(new_n224), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n229), .A2(new_n244), .A3(new_n231), .A4(new_n239), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n215), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT67), .B1(new_n237), .B2(G131), .ZN(new_n247));
  AOI211_X1 g061(.A(new_n232), .B(new_n230), .C1(new_n235), .C2(new_n236), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n231), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n226), .A2(new_n228), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT69), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n246), .A2(KEYINPUT70), .A3(new_n224), .A4(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n224), .A3(new_n215), .A4(new_n245), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n245), .A3(new_n215), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n252), .A2(new_n255), .B1(new_n223), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n243), .B1(new_n257), .B2(new_n242), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n260), .B(KEYINPUT27), .Z(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n187), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n252), .A2(new_n255), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n215), .A2(new_n270), .A3(new_n240), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n256), .B2(KEYINPUT30), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n224), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n263), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n252), .A2(new_n255), .A3(KEYINPUT28), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n224), .B1(new_n215), .B2(new_n240), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n241), .B2(new_n242), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n274), .B(new_n275), .C1(new_n263), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n268), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n266), .A2(new_n267), .ZN(new_n282));
  OAI21_X1  g096(.A(G472), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n269), .B(new_n264), .C1(new_n224), .C2(new_n272), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n215), .A2(new_n245), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n289), .A2(new_n230), .B1(new_n234), .B2(new_n238), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n244), .B1(new_n290), .B2(new_n229), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT30), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n215), .A2(new_n270), .A3(new_n240), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n223), .B1(new_n252), .B2(new_n255), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n287), .B1(new_n295), .B2(new_n264), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n284), .B1(new_n286), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n279), .A2(new_n263), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n263), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n284), .B1(new_n285), .B2(KEYINPUT31), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n297), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n283), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G234), .ZN(new_n312));
  OAI21_X1  g126(.A(G217), .B1(new_n312), .B2(G902), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT74), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OR3_X1    g129(.A1(new_n227), .A2(KEYINPUT75), .A3(G119), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n316), .B(new_n319), .C1(new_n317), .C2(G128), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT24), .B(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n317), .A2(G128), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n318), .B(new_n323), .C1(new_n324), .C2(KEYINPUT23), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(G110), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT76), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G146), .ZN(new_n336));
  XNOR2_X1  g150(.A(G125), .B(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n192), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n326), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n331), .A2(new_n192), .A3(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n325), .A2(G110), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n341), .B(new_n342), .C1(new_n321), .C2(new_n320), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT22), .B(G137), .ZN(new_n345));
  INV_X1    g159(.A(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n339), .A2(new_n343), .A3(new_n348), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n187), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(KEYINPUT78), .B2(KEYINPUT25), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n350), .A2(KEYINPUT77), .A3(new_n187), .A4(new_n351), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n357), .A2(KEYINPUT78), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n315), .B(new_n356), .C1(new_n358), .C2(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n313), .A2(new_n187), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT79), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n350), .A2(new_n361), .A3(new_n351), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n311), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  OAI21_X1  g180(.A(G221), .B1(new_n366), .B2(G902), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n367), .B(KEYINPUT80), .Z(new_n368));
  INV_X1    g182(.A(G469), .ZN(new_n369));
  INV_X1    g183(.A(new_n213), .ZN(new_n370));
  INV_X1    g184(.A(new_n214), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT83), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G104), .B(G107), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G104), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G107), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G101), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n376), .A3(G104), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n383), .A2(new_n385), .A3(new_n374), .A4(new_n379), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n375), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n250), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n387), .A2(new_n250), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n372), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT12), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n372), .B(KEYINPUT12), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n383), .A2(new_n385), .A3(new_n379), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n399), .A2(new_n200), .B1(new_n388), .B2(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n370), .A2(new_n371), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n388), .B2(KEYINPUT10), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT10), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT82), .B(new_n405), .C1(new_n387), .C2(new_n250), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n400), .A2(new_n402), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G140), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n346), .A2(G227), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n394), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT85), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n399), .A2(new_n200), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n388), .A2(KEYINPUT10), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n414), .A2(new_n404), .A3(new_n415), .A4(new_n406), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(KEYINPUT84), .B2(new_n402), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n402), .A2(KEYINPUT84), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(new_n400), .A3(new_n404), .A4(new_n406), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n410), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT86), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n422), .A3(new_n410), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n369), .B(new_n187), .C1(new_n413), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n410), .B1(new_n417), .B2(new_n419), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n411), .B1(new_n394), .B2(new_n407), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G469), .B1(new_n428), .B2(G902), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n368), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(G143), .B1(new_n259), .B2(G214), .ZN(new_n433));
  OAI21_X1  g247(.A(G131), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n230), .A3(new_n431), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(KEYINPUT17), .B(G131), .C1(new_n432), .C2(new_n433), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n438), .A2(new_n336), .A3(new_n340), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT18), .A2(G131), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n431), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n338), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT18), .B(G131), .C1(new_n432), .C2(new_n433), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(G113), .B(G122), .Z(new_n448));
  XOR2_X1   g262(.A(KEYINPUT91), .B(G104), .Z(new_n449));
  XOR2_X1   g263(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT90), .B1(new_n337), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n329), .A2(KEYINPUT19), .A3(new_n330), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n329), .A2(KEYINPUT90), .A3(KEYINPUT19), .A4(new_n330), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n192), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n434), .A2(new_n436), .B1(G146), .B2(new_n335), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n458), .A2(new_n459), .B1(new_n446), .B2(new_n445), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n451), .B1(new_n460), .B2(new_n450), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n462));
  NOR2_X1   g276(.A1(G475), .A2(G902), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n463), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n447), .ZN(new_n467));
  INV_X1    g281(.A(new_n450), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n469), .B2(new_n451), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n471));
  OAI21_X1  g285(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n451), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n450), .B1(new_n440), .B2(new_n447), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n187), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(G234), .A2(G237), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n478), .A2(G952), .A3(new_n346), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n478), .A2(G902), .A3(G953), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(G898), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G128), .B(G143), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT13), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n194), .A2(G128), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n484), .B(G134), .C1(KEYINPUT13), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n227), .A2(G143), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n483), .A2(KEYINPUT93), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n493));
  INV_X1    g307(.A(G122), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(G116), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G116), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n496), .A2(KEYINPUT92), .A3(G122), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n495), .A2(new_n497), .B1(G116), .B2(new_n494), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n498), .A2(G107), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(G107), .ZN(new_n500));
  OAI221_X1 g314(.A(new_n486), .B1(new_n492), .B2(G134), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n495), .B2(new_n497), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n502), .A3(G107), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n490), .A2(new_n491), .A3(G134), .ZN(new_n505));
  AOI21_X1  g319(.A(G134), .B1(new_n490), .B2(new_n491), .ZN(new_n506));
  OAI221_X1 g320(.A(new_n503), .B1(new_n498), .B2(new_n504), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G217), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n366), .A2(new_n508), .A3(G953), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n501), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n501), .B2(new_n507), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n187), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G478), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI221_X1 g329(.A(new_n187), .B1(KEYINPUT15), .B2(new_n513), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n477), .A2(new_n482), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n221), .A2(new_n222), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n222), .A2(KEYINPUT5), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n496), .A2(G119), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n218), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n387), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n398), .A2(new_n396), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n223), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G122), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(new_n530), .A3(new_n532), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT6), .A3(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n200), .A2(new_n333), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n250), .A2(new_n333), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n346), .A2(G224), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT87), .Z(new_n540));
  AND3_X1   g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n537), .B2(new_n538), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n531), .A2(new_n544), .A3(new_n533), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n536), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n537), .A2(KEYINPUT7), .A3(new_n538), .A4(new_n539), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n548));
  AOI21_X1  g362(.A(G125), .B1(new_n226), .B2(new_n228), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n550));
  OAI22_X1  g364(.A1(new_n200), .A2(new_n333), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n538), .A2(KEYINPUT88), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n532), .B(KEYINPUT8), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n525), .A2(new_n387), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n526), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n535), .A2(new_n547), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n557), .A2(new_n187), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n546), .B2(new_n558), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G214), .B1(G237), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n430), .A2(new_n518), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n365), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n374), .ZN(G3));
  INV_X1    g383(.A(new_n482), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n570), .B(new_n564), .C1(new_n561), .C2(new_n562), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n363), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n430), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n305), .A2(new_n187), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n574), .A2(G472), .B1(new_n307), .B2(new_n305), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n510), .A2(new_n511), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT33), .B1(new_n511), .B2(KEYINPUT94), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G478), .ZN(new_n583));
  MUX2_X1   g397(.A(new_n187), .B(new_n512), .S(new_n513), .Z(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n477), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT34), .B(G104), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  XNOR2_X1  g403(.A(new_n470), .B(new_n471), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n590), .A2(new_n476), .A3(new_n517), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n576), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G107), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G9));
  OAI21_X1  g410(.A(new_n344), .B1(KEYINPUT36), .B2(new_n349), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n339), .A2(new_n343), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n361), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT97), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n359), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n356), .A2(new_n315), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT25), .B1(new_n357), .B2(KEYINPUT78), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n600), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT98), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n430), .A2(new_n566), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n518), .A3(new_n575), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT37), .B(G110), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G12));
  INV_X1    g428(.A(G900), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n479), .B1(new_n480), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n590), .A2(new_n517), .A3(new_n476), .A4(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n311), .A2(new_n611), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G128), .ZN(G30));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  OR3_X1    g436(.A1(new_n257), .A2(KEYINPUT99), .A3(new_n264), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT99), .B1(new_n257), .B2(new_n264), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n285), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(new_n187), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n309), .A2(new_n310), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n563), .B(KEYINPUT38), .Z(new_n628));
  NOR2_X1   g442(.A1(new_n606), .A2(new_n608), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n472), .A2(new_n476), .B1(new_n515), .B2(new_n516), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n630), .A2(new_n565), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n634), .A2(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(KEYINPUT100), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n616), .B(KEYINPUT39), .Z(new_n637));
  NAND2_X1  g451(.A1(new_n430), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT40), .Z(new_n639));
  NAND3_X1  g453(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G143), .ZN(G45));
  NOR2_X1   g455(.A1(new_n585), .A2(new_n616), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n311), .A2(new_n611), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  OAI21_X1  g458(.A(new_n187), .B1(new_n413), .B2(new_n424), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G469), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n646), .A2(new_n425), .ZN(new_n647));
  INV_X1    g461(.A(new_n368), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n585), .A2(new_n571), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n649), .A2(new_n311), .A3(new_n364), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  AND3_X1   g467(.A1(new_n566), .A2(new_n570), .A3(new_n591), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n649), .A2(new_n311), .A3(new_n364), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G116), .ZN(G18));
  NAND4_X1  g470(.A1(new_n646), .A2(new_n566), .A3(new_n648), .A4(new_n425), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n610), .A2(new_n518), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n311), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G119), .ZN(G21));
  AOI21_X1  g475(.A(new_n622), .B1(new_n305), .B2(new_n187), .ZN(new_n662));
  INV_X1    g476(.A(new_n307), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n295), .A2(new_n287), .A3(new_n264), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n258), .A2(new_n263), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n662), .A2(new_n363), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n631), .B(new_n564), .C1(new_n561), .C2(new_n562), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n482), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n648), .A2(new_n672), .A3(new_n425), .A4(new_n646), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT101), .B(G122), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G24));
  NAND4_X1  g490(.A1(new_n647), .A2(new_n566), .A3(new_n648), .A4(new_n642), .ZN(new_n677));
  INV_X1    g491(.A(new_n669), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n303), .B1(new_n666), .B2(new_n284), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(new_n302), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n630), .B(new_n678), .C1(new_n680), .C2(new_n622), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n574), .A2(G472), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(KEYINPUT102), .A3(new_n630), .A4(new_n678), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n677), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n333), .ZN(G27));
  NAND2_X1  g501(.A1(new_n546), .A2(new_n558), .ZN(new_n688));
  INV_X1    g502(.A(new_n559), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n564), .A3(new_n560), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT103), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n642), .A2(new_n692), .A3(new_n430), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n311), .A3(new_n364), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT104), .B(G131), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G33));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n618), .B(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n692), .A2(new_n701), .A3(new_n430), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n311), .A2(new_n702), .A3(new_n364), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G134), .ZN(G36));
  NAND2_X1  g518(.A1(new_n583), .A2(new_n584), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(new_n477), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT43), .Z(new_n707));
  OR2_X1    g521(.A1(new_n575), .A2(new_n629), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n428), .A2(KEYINPUT45), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n428), .A2(KEYINPUT45), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(G469), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(G469), .A2(G902), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT46), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(KEYINPUT46), .A3(new_n720), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n425), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n368), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n637), .A3(new_n692), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n715), .A2(new_n716), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G137), .ZN(G39));
  XNOR2_X1  g544(.A(new_n727), .B(KEYINPUT47), .ZN(new_n731));
  INV_X1    g545(.A(new_n692), .ZN(new_n732));
  INV_X1    g546(.A(new_n642), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n311), .A2(new_n732), .A3(new_n364), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  NOR2_X1   g550(.A1(new_n626), .A2(new_n622), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n305), .A2(new_n307), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT32), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n737), .B1(new_n739), .B2(new_n308), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n364), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n647), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n647), .A2(new_n743), .ZN(new_n745));
  NOR4_X1   g559(.A1(new_n628), .A2(new_n706), .A3(new_n565), .A4(new_n368), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n742), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT113), .B1(new_n649), .B2(new_n692), .ZN(new_n748));
  INV_X1    g562(.A(new_n479), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n649), .A2(KEYINPUT113), .A3(new_n692), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n707), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT114), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n683), .A2(new_n685), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n707), .A2(new_n479), .A3(new_n670), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n647), .A2(new_n368), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n692), .B(new_n757), .C1(new_n731), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n628), .A2(new_n564), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n649), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n756), .A2(new_n760), .A3(new_n762), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n750), .A2(new_n751), .A3(new_n742), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n477), .B1(new_n583), .B2(new_n584), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n755), .A2(new_n759), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n755), .A2(KEYINPUT51), .A3(new_n759), .A4(new_n767), .ZN(new_n771));
  INV_X1    g585(.A(new_n365), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n753), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT48), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n753), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(G952), .B(new_n346), .C1(new_n756), .C2(new_n657), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n765), .B2(new_n586), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n770), .A2(new_n771), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n733), .A2(new_n657), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n669), .B1(new_n574), .B2(G472), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT102), .B1(new_n782), .B2(new_n630), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n662), .A2(new_n682), .A3(new_n629), .A4(new_n669), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n620), .A3(new_n643), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n630), .A2(new_n616), .A3(new_n632), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n430), .A3(new_n566), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n740), .A2(KEYINPUT111), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n790));
  INV_X1    g604(.A(new_n788), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n627), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n620), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n686), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT111), .B1(new_n740), .B2(new_n788), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n627), .A2(new_n790), .A3(new_n791), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n797), .A3(new_n643), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n651), .A2(new_n655), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n517), .B(KEYINPUT108), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n585), .B1(new_n477), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n573), .A2(new_n575), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n660), .A2(new_n612), .A3(new_n674), .A4(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n802), .A2(new_n806), .A3(new_n568), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n794), .A2(new_n801), .A3(new_n807), .A4(new_n697), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n590), .A2(new_n476), .A3(new_n617), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n803), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n430), .A2(new_n692), .A3(new_n610), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n311), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n703), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT109), .B1(new_n754), .B2(new_n694), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n818), .B(new_n693), .C1(new_n683), .C2(new_n685), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT110), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n694), .B1(new_n783), .B2(new_n784), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n754), .A2(KEYINPUT109), .A3(new_n694), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n816), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n809), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n825), .B2(new_n816), .ZN(new_n830));
  AOI211_X1 g644(.A(KEYINPUT110), .B(new_n815), .C1(new_n823), .C2(new_n824), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n795), .B2(new_n686), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n832), .A2(new_n808), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n834), .B1(new_n832), .B2(new_n808), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n794), .A2(new_n697), .A3(new_n807), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n828), .A3(new_n801), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n840), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n839), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n840), .A2(new_n845), .A3(new_n844), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n841), .A2(new_n828), .A3(new_n801), .A4(new_n835), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n780), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  INV_X1    g667(.A(G952), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n346), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n747), .B1(new_n856), .B2(new_n857), .ZN(G75));
  NOR2_X1   g672(.A1(new_n346), .A2(G952), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n840), .A2(new_n844), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n861), .A2(G210), .A3(G902), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n536), .A2(new_n545), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(new_n543), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n860), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n187), .B1(new_n840), .B2(new_n844), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n871), .A2(new_n869), .A3(G210), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n865), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT117), .B(new_n865), .C1(new_n870), .C2(new_n872), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(G51));
  INV_X1    g691(.A(new_n719), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(KEYINPUT118), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n413), .A2(new_n424), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n832), .A2(new_n808), .A3(new_n842), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(new_n829), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n846), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n720), .B(KEYINPUT57), .Z(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n860), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT119), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n892), .B(new_n860), .C1(new_n883), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  INV_X1    g709(.A(new_n461), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n859), .ZN(G60));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n513), .A2(new_n187), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT59), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n582), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT120), .B1(new_n887), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  INV_X1    g719(.A(new_n903), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n905), .B(new_n906), .C1(new_n886), .C2(new_n846), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n860), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n851), .A2(new_n847), .ZN(new_n909));
  INV_X1    g723(.A(new_n902), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n581), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n900), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n848), .A2(new_n850), .A3(KEYINPUT112), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n839), .B1(new_n838), .B2(new_n846), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n582), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n845), .B1(new_n840), .B2(new_n844), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n903), .B1(new_n848), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n903), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n859), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(KEYINPUT121), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n912), .A2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  AND2_X1   g739(.A1(new_n861), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n597), .A2(new_n599), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n860), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n861), .A2(new_n925), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n350), .A2(new_n351), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G66));
  INV_X1    g752(.A(G224), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n481), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n807), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n863), .B1(G898), .B2(new_n346), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  AND2_X1   g758(.A1(new_n735), .A2(new_n697), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n786), .B(KEYINPUT125), .Z(new_n946));
  AND4_X1   g760(.A1(new_n566), .A2(new_n727), .A3(new_n631), .A4(new_n637), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n772), .B1(new_n947), .B2(new_n702), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n945), .A2(new_n729), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n294), .B(new_n457), .ZN(new_n951));
  NAND2_X1  g765(.A1(G900), .A2(G953), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n804), .B(KEYINPUT126), .Z(new_n955));
  OR4_X1    g769(.A1(new_n365), .A2(new_n955), .A3(new_n638), .A4(new_n732), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n729), .A2(new_n735), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n946), .A2(new_n640), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n954), .B1(new_n963), .B2(new_n951), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n346), .B1(G227), .B2(G900), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n965), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n954), .B(new_n967), .C1(new_n963), .C2(new_n951), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(new_n962), .A2(new_n807), .ZN(new_n970));
  XNOR2_X1  g784(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n263), .B(new_n295), .C1(new_n970), .C2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n807), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n949), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n263), .A3(new_n295), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n860), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n274), .A2(new_n285), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n973), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n840), .B2(new_n849), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(G57));
endmodule


