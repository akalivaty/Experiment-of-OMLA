//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  OR2_X1    g0003(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n205));
  NAND3_X1  g0005(.A1(new_n204), .A2(G50), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g0006(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n206), .A2(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n216), .B(new_n222), .C1(G97), .C2(G257), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G1), .B2(G20), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  AOI211_X1 g0025(.A(new_n212), .B(new_n225), .C1(new_n211), .C2(new_n210), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  AND2_X1   g0041(.A1(KEYINPUT3), .A2(G33), .ZN(new_n242));
  NOR2_X1   g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G20), .ZN(new_n245));
  AOI21_X1  g0045(.A(KEYINPUT7), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT7), .ZN(new_n247));
  NOR4_X1   g0047(.A1(new_n242), .A2(new_n243), .A3(new_n247), .A4(G20), .ZN(new_n248));
  OAI21_X1  g0048(.A(G68), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G159), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G58), .A2(G68), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT75), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n254), .B2(new_n203), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT16), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n249), .A2(KEYINPUT16), .A3(new_n251), .A4(new_n255), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT66), .B(G1), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT70), .ZN(new_n265));
  INV_X1    g0065(.A(G13), .ZN(new_n266));
  NOR4_X1   g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .A4(new_n245), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n245), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT70), .B1(new_n272), .B2(G13), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  INV_X1    g0075(.A(G58), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT8), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT8), .B(G58), .Z(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n270), .A2(G1), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n282));
  OAI211_X1 g0082(.A(G13), .B(G20), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n265), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n272), .A2(KEYINPUT70), .A3(G13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n261), .ZN(new_n287));
  INV_X1    g0087(.A(new_n272), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n289), .A2(new_n279), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n263), .A2(new_n280), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G41), .A2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n294), .A2(new_n268), .A3(G274), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT67), .B1(new_n264), .B2(new_n293), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n269), .A2(new_n271), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(new_n294), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n295), .B1(new_n303), .B2(G232), .ZN(new_n304));
  OR2_X1    g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G223), .B2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(G1698), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G226), .ZN(new_n310));
  INV_X1    g0110(.A(G33), .ZN(new_n311));
  INV_X1    g0111(.A(G87), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n308), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n298), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n304), .A2(G190), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n304), .B2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n292), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT17), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n292), .A2(KEYINPUT17), .A3(new_n315), .A4(new_n318), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n304), .A2(new_n324), .A3(new_n314), .ZN(new_n325));
  AOI21_X1  g0125(.A(G169), .B1(new_n304), .B2(new_n314), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n291), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT18), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT18), .B1(new_n291), .B2(new_n327), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n335), .A2(KEYINPUT76), .A3(KEYINPUT77), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n330), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n333), .A3(new_n331), .ZN(new_n338));
  INV_X1    g0138(.A(new_n330), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT77), .B1(new_n335), .B2(KEYINPUT76), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n323), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT65), .B(G226), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n295), .B1(new_n303), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n244), .B1(G222), .B2(new_n309), .ZN(new_n345));
  INV_X1    g0145(.A(G223), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n309), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G77), .B2(new_n307), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(new_n297), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n245), .A2(G33), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT69), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G150), .ZN(new_n355));
  INV_X1    g0155(.A(new_n250), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n279), .A2(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n245), .B1(new_n203), .B2(new_n218), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n261), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n274), .A2(new_n218), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n218), .C2(new_n289), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n351), .B(new_n361), .C1(G179), .C2(new_n349), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT71), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n356), .A2(new_n218), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n245), .A2(G68), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n352), .B(KEYINPUT69), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(G77), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT11), .B1(new_n368), .B2(new_n287), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT11), .ZN(new_n370));
  INV_X1    g0170(.A(G77), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n354), .A2(new_n371), .B1(new_n245), .B2(G68), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n261), .C1(new_n372), .C2(new_n365), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n289), .A2(new_n220), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT12), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n274), .A2(new_n376), .A3(new_n220), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT12), .B1(new_n286), .B2(G68), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n295), .B1(new_n303), .B2(G238), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n307), .B1(G232), .B2(new_n309), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G226), .A2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n298), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT13), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n381), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n380), .B1(new_n391), .B2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n381), .B2(new_n386), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G190), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n295), .B1(new_n303), .B2(G244), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n244), .B1(G232), .B2(new_n309), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n221), .B2(new_n309), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G107), .B2(new_n307), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n297), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n402), .A2(G179), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n278), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n406), .A2(new_n352), .B1(new_n356), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n245), .A2(new_n371), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n261), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n274), .A2(new_n371), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n371), .C2(new_n289), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n402), .A2(new_n350), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n403), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n364), .A2(new_n397), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n380), .B(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(G169), .B1(new_n393), .B2(new_n394), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n391), .A2(new_n420), .A3(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n395), .A2(G179), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n415), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT9), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n361), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G190), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n349), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n361), .A2(new_n425), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n349), .A2(G200), .B1(KEYINPUT73), .B2(KEYINPUT10), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n426), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(KEYINPUT73), .A2(KEYINPUT10), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n412), .B1(G200), .B2(new_n402), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n402), .A2(new_n427), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n342), .A2(new_n424), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G97), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n274), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n264), .A2(new_n311), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n286), .A2(G97), .A3(new_n287), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n305), .A2(new_n245), .A3(new_n306), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n247), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n244), .A2(KEYINPUT7), .A3(new_n245), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n250), .A2(G77), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT6), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n440), .A2(new_n445), .ZN(new_n453));
  NOR2_X1   g0253(.A1(G97), .A2(G107), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n445), .A2(KEYINPUT6), .A3(G97), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n245), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n449), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n441), .B(new_n444), .C1(new_n458), .C2(new_n287), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT79), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(G107), .B1(new_n246), .B2(new_n248), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n455), .A2(new_n456), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n450), .C1(new_n245), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n261), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n465), .A2(KEYINPUT79), .A3(new_n441), .A4(new_n444), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n307), .A2(G250), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n309), .B1(new_n468), .B2(KEYINPUT4), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1698), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(G244), .C1(new_n243), .C2(new_n242), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  INV_X1    g0273(.A(G244), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n305), .B2(new_n306), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n472), .B(new_n473), .C1(new_n475), .C2(KEYINPUT4), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n298), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G45), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n269), .B2(new_n271), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT5), .B(G41), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(G274), .A3(new_n297), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n298), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT78), .A3(G257), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT78), .B1(new_n482), .B2(G257), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n477), .B(new_n481), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G169), .ZN(new_n487));
  INV_X1    g0287(.A(new_n485), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n483), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(G179), .A3(new_n481), .A4(new_n477), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n467), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n459), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n486), .A2(G200), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n427), .C2(new_n486), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n221), .A2(new_n309), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n474), .A2(G1698), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n498), .C1(new_n242), .C2(new_n243), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G116), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n297), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n300), .A2(G45), .A3(G274), .A4(new_n297), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT80), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n479), .A2(new_n504), .A3(G274), .A4(new_n297), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G250), .B(new_n297), .C1(new_n264), .C2(new_n478), .ZN(new_n507));
  AOI21_X1  g0307(.A(G169), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(new_n501), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n509), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n324), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT19), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n245), .B1(new_n382), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n312), .A2(new_n440), .A3(new_n445), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT81), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n307), .A2(new_n245), .A3(G68), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n520), .A3(new_n516), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n514), .B1(new_n352), .B2(new_n440), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n274), .A2(new_n406), .B1(new_n523), .B2(new_n261), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n404), .B(KEYINPUT72), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n286), .A2(new_n287), .A3(new_n525), .A4(new_n443), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n513), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n274), .A2(new_n406), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n261), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n513), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n512), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n506), .A2(G190), .A3(new_n507), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n286), .A2(G87), .A3(new_n287), .A4(new_n443), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n524), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n509), .A2(new_n507), .A3(new_n510), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n496), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G257), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G1698), .ZN(new_n541));
  OAI221_X1 g0341(.A(new_n541), .B1(G250), .B2(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n298), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n482), .A2(G264), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n427), .A4(new_n481), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT88), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT87), .ZN(new_n549));
  INV_X1    g0349(.A(G264), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n550), .B(new_n298), .C1(new_n479), .C2(new_n480), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n297), .B1(new_n542), .B2(new_n543), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT87), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n481), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n316), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n261), .B(new_n442), .C1(new_n284), .C2(new_n285), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G107), .ZN(new_n559));
  AND2_X1   g0359(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n560));
  NOR2_X1   g0360(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n307), .A2(new_n562), .A3(new_n245), .A4(G87), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n245), .B(G87), .C1(new_n242), .C2(new_n243), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n445), .A2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n245), .A2(G33), .A3(G116), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n563), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n571), .B(new_n572), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n573), .A2(new_n287), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n445), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n286), .B2(G107), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n557), .A2(new_n559), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n559), .B(new_n578), .C1(new_n573), .C2(new_n287), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n545), .A2(new_n546), .A3(new_n481), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n555), .B2(new_n324), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n284), .A2(new_n214), .A3(new_n285), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n214), .A2(G20), .ZN(new_n588));
  AOI21_X1  g0388(.A(G20), .B1(G33), .B2(G283), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n311), .A2(G97), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT85), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT85), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n261), .B(new_n588), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n587), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT84), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n287), .B(new_n443), .C1(new_n267), .C2(new_n273), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n214), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n558), .A2(KEYINPUT84), .A3(G116), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n540), .A2(G1698), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n550), .A2(new_n309), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n307), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G303), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n307), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n605), .B(KEYINPUT83), .C1(new_n606), .C2(new_n307), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n298), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n482), .A2(G270), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n481), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G169), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n586), .B1(new_n602), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(G200), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n602), .B(new_n617), .C1(new_n427), .C2(new_n614), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n593), .A2(new_n594), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n593), .A2(new_n594), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n619), .A2(new_n620), .B1(new_n214), .B2(new_n274), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT84), .B1(new_n558), .B2(G116), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n599), .A2(new_n598), .A3(new_n214), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n350), .B1(new_n611), .B2(new_n613), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(KEYINPUT21), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n614), .A2(new_n324), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n616), .A2(new_n618), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n439), .A2(new_n539), .A3(new_n585), .A4(new_n629), .ZN(G372));
  NAND2_X1  g0430(.A1(new_n423), .A2(new_n417), .ZN(new_n631));
  INV_X1    g0431(.A(new_n397), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n414), .ZN(new_n633));
  INV_X1    g0433(.A(new_n323), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n339), .B2(new_n332), .ZN(new_n635));
  INV_X1    g0435(.A(new_n433), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n364), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n506), .A2(new_n324), .A3(new_n507), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n511), .B2(G169), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n524), .A2(new_n513), .A3(new_n526), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT82), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n524), .A2(new_n532), .A3(new_n533), .ZN(new_n645));
  AOI211_X1 g0445(.A(KEYINPUT89), .B(new_n316), .C1(new_n506), .C2(new_n507), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n535), .B2(G200), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT90), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n648), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n535), .A2(new_n647), .A3(G200), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n534), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n531), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n491), .A2(new_n459), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT26), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n461), .A2(new_n466), .B1(new_n487), .B2(new_n490), .ZN(new_n660));
  XOR2_X1   g0460(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n537), .A3(new_n531), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT92), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n645), .B1(G200), .B2(new_n535), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n644), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT92), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n660), .A4(new_n661), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n494), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n486), .A2(new_n427), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n670), .A2(new_n671), .A3(new_n459), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n660), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n531), .A2(new_n653), .A3(new_n654), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n654), .B1(new_n531), .B2(new_n653), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n616), .A2(new_n626), .A3(new_n584), .A4(new_n628), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n579), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n531), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n669), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n638), .B1(new_n438), .B2(new_n680), .ZN(G369));
  NAND2_X1  g0481(.A1(new_n245), .A2(G13), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n264), .A2(KEYINPUT27), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT27), .B1(new_n264), .B2(new_n682), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G213), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n602), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n629), .A2(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n629), .A2(KEYINPUT93), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n616), .A2(new_n626), .A3(new_n628), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT94), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n580), .A2(new_n687), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n585), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n584), .B2(new_n688), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n677), .A2(new_n579), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n688), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n209), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n516), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n206), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n661), .B1(new_n665), .B2(new_n660), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n657), .B1(new_n650), .B2(new_n655), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(KEYINPUT26), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n688), .B1(new_n679), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n688), .B1(new_n669), .B2(new_n679), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(KEYINPUT29), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n539), .A2(new_n585), .A3(new_n629), .A4(new_n688), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n553), .A2(new_n554), .ZN(new_n721));
  INV_X1    g0521(.A(new_n486), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n627), .A2(new_n721), .A3(new_n511), .A4(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n511), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n486), .A3(new_n614), .A4(new_n555), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n724), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n687), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n720), .A2(new_n730), .A3(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n732), .A3(new_n687), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(G330), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n719), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n712), .B1(new_n736), .B2(G1), .ZN(G364));
  XNOR2_X1  g0537(.A(new_n682), .B(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G1), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n707), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n324), .A2(new_n316), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n245), .A2(new_n427), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n245), .A2(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n324), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G50), .A2(new_n746), .B1(new_n750), .B2(G77), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(new_n748), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n276), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n743), .A2(new_n747), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n755), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n753), .B1(G68), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n747), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  OR3_X1    g0564(.A1(new_n763), .A2(KEYINPUT32), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(KEYINPUT32), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n316), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n747), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n765), .B(new_n766), .C1(new_n445), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n245), .B1(new_n762), .B2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n440), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n769), .A2(new_n244), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n744), .A2(new_n767), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n761), .B(new_n772), .C1(new_n312), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n244), .B1(new_n773), .B2(new_n606), .ZN(new_n776));
  INV_X1    g0576(.A(new_n752), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G322), .A2(new_n777), .B1(new_n750), .B2(G311), .ZN(new_n778));
  INV_X1    g0578(.A(G329), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n779), .B2(new_n763), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n776), .B(new_n780), .C1(new_n760), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n745), .A2(new_n783), .B1(new_n770), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT98), .Z(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n782), .B(new_n786), .C1(new_n787), .C2(new_n768), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n260), .B1(G20), .B2(new_n350), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n742), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n791), .B1(new_n697), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(new_n790), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n237), .A2(G45), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n706), .A2(new_n307), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G45), .C2(new_n206), .ZN(new_n800));
  INV_X1    g0600(.A(G355), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n307), .A2(new_n209), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(G116), .B2(new_n209), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n796), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT99), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n698), .A2(new_n741), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G330), .B2(new_n697), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NOR2_X1   g0609(.A1(new_n414), .A2(new_n687), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n434), .A2(new_n435), .B1(new_n412), .B2(new_n687), .ZN(new_n812));
  INV_X1    g0612(.A(new_n414), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n718), .B(new_n815), .ZN(new_n816));
  OR3_X1    g0616(.A1(new_n816), .A2(new_n735), .A3(KEYINPUT102), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT102), .B1(new_n816), .B2(new_n735), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n735), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n817), .A2(new_n742), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G137), .A2(new_n746), .B1(new_n777), .B2(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n764), .B2(new_n749), .C1(new_n759), .C2(new_n355), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT34), .ZN(new_n823));
  INV_X1    g0623(.A(new_n768), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G68), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n307), .B1(new_n763), .B2(new_n826), .C1(new_n218), .C2(new_n773), .ZN(new_n827));
  INV_X1    g0627(.A(new_n770), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(G58), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n823), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n244), .B1(new_n763), .B2(new_n831), .C1(new_n312), .C2(new_n768), .ZN(new_n832));
  INV_X1    g0632(.A(new_n773), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n771), .B(new_n832), .C1(G107), .C2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n752), .A2(new_n784), .B1(new_n749), .B2(new_n214), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n760), .B2(G283), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n606), .C2(new_n745), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT101), .Z(new_n839));
  AOI21_X1  g0639(.A(new_n742), .B1(new_n839), .B2(new_n790), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n790), .A2(new_n792), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n371), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n840), .B(new_n843), .C1(new_n793), .C2(new_n815), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n820), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  AOI22_X1  g0646(.A1(new_n417), .A2(new_n687), .B1(new_n392), .B2(new_n396), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n423), .A2(new_n417), .A3(KEYINPUT104), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT104), .B1(new_n423), .B2(new_n417), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n417), .B(new_n687), .C1(new_n632), .C2(new_n423), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n852), .A2(new_n731), .A3(new_n733), .A4(new_n815), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n634), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n685), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n291), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n291), .B1(new_n327), .B2(new_n858), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n319), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n319), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n869), .B(new_n866), .C1(new_n857), .C2(new_n860), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n854), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(KEYINPUT38), .B(new_n867), .C1(new_n342), .C2(new_n859), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n339), .A2(new_n332), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n859), .B1(new_n634), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n869), .B1(new_n876), .B2(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n854), .A3(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n731), .A2(new_n733), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n438), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(G330), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n815), .B(new_n688), .C1(new_n669), .C2(new_n679), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n885), .A2(KEYINPUT103), .A3(new_n811), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT103), .B1(new_n885), .B2(new_n811), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n852), .B1(new_n868), .B2(new_n870), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n867), .B1(new_n342), .B2(new_n859), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n869), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n878), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n848), .A2(new_n849), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n688), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n339), .A2(new_n332), .A3(new_n685), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n637), .B1(new_n719), .B2(new_n439), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n884), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n300), .B2(new_n738), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT35), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n207), .B1(new_n463), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(G116), .C1(new_n904), .C2(new_n463), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n254), .A2(new_n371), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n908), .A2(new_n206), .B1(G50), .B2(new_n220), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n266), .A3(new_n264), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(G367));
  OAI21_X1  g0711(.A(new_n244), .B1(new_n768), .B2(new_n440), .ZN(new_n912));
  INV_X1    g0712(.A(new_n763), .ZN(new_n913));
  AOI22_X1  g0713(.A1(G283), .A2(new_n750), .B1(new_n913), .B2(G317), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n914), .B1(new_n606), .B2(new_n752), .C1(new_n831), .C2(new_n745), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n912), .B(new_n915), .C1(G107), .C2(new_n828), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n833), .A2(G116), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT46), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n916), .B(new_n918), .C1(new_n784), .C2(new_n759), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT109), .ZN(new_n920));
  INV_X1    g0720(.A(G143), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n745), .A2(new_n921), .B1(new_n752), .B2(new_n355), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n760), .B2(G159), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n307), .B1(new_n773), .B2(new_n276), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n768), .A2(new_n371), .B1(new_n770), .B2(new_n220), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n924), .B(new_n925), .C1(G137), .C2(new_n913), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n923), .B(new_n926), .C1(new_n218), .C2(new_n749), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT110), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT47), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n742), .B1(new_n930), .B2(new_n790), .ZN(new_n931));
  INV_X1    g0731(.A(new_n799), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n797), .B1(new_n406), .B2(new_n209), .C1(new_n233), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n524), .A2(new_n533), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n687), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n656), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n531), .B2(new_n935), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n931), .B(new_n933), .C1(new_n795), .C2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n740), .B(KEYINPUT108), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n698), .A2(new_n701), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n673), .B1(new_n493), .B2(new_n688), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n658), .A2(new_n687), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n704), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT45), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n704), .A2(new_n673), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT106), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n693), .A2(new_n688), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n585), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n701), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n952), .A2(new_n955), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n736), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n702), .B(new_n949), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n736), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n707), .B(KEYINPUT41), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n940), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n941), .A2(new_n944), .ZN(new_n964));
  INV_X1    g0764(.A(new_n944), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n492), .B1(new_n965), .B2(new_n584), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT105), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n688), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n954), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT42), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n937), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n964), .B(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n938), .B1(new_n963), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT111), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n977), .B(new_n938), .C1(new_n963), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(G387));
  NAND2_X1  g0779(.A1(new_n957), .A2(new_n956), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n735), .B2(new_n719), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n957), .A2(new_n736), .A3(new_n956), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n707), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n957), .A2(new_n956), .A3(new_n940), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n745), .A2(new_n764), .B1(new_n749), .B2(new_n220), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n307), .B1(new_n768), .B2(new_n440), .C1(new_n218), .C2(new_n752), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G150), .C2(new_n913), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n833), .A2(G77), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n759), .A2(new_n279), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n525), .A2(new_n828), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G322), .A2(new_n746), .B1(new_n777), .B2(G317), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n606), .B2(new_n749), .C1(new_n759), .C2(new_n831), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n787), .B2(new_n770), .C1(new_n784), .C2(new_n773), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT49), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n244), .B1(new_n763), .B2(new_n783), .C1(new_n214), .C2(new_n768), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT112), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n991), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n799), .B1(new_n230), .B2(new_n478), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n709), .B2(new_n802), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n220), .A2(new_n371), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n278), .A2(new_n218), .ZN(new_n1003));
  AOI211_X1 g0803(.A(G116), .B(new_n516), .C1(new_n1003), .C2(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n478), .C1(KEYINPUT50), .C2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1001), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(G107), .B2(new_n209), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n999), .A2(new_n790), .B1(new_n797), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n741), .C1(new_n701), .C2(new_n795), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n984), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n983), .A2(new_n1010), .ZN(G393));
  INV_X1    g0811(.A(new_n982), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n707), .B1(new_n1012), .B2(new_n959), .C1(new_n960), .C2(new_n958), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n797), .B1(new_n440), .B2(new_n209), .C1(new_n240), .C2(new_n932), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n944), .A2(new_n795), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT113), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G68), .A2(new_n833), .B1(new_n913), .B2(G143), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n371), .B2(new_n770), .C1(new_n407), .C2(new_n749), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n307), .B1(new_n768), .B2(new_n312), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n745), .A2(new_n355), .B1(new_n752), .B2(new_n764), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n218), .C2(new_n759), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G294), .A2(new_n750), .B1(new_n913), .B2(G322), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n445), .B2(new_n768), .C1(new_n787), .C2(new_n773), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n307), .B(new_n1026), .C1(G116), .C2(new_n828), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n606), .B2(new_n759), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G317), .A2(new_n746), .B1(new_n777), .B2(G311), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT52), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1024), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n742), .B1(new_n1031), .B2(new_n790), .ZN(new_n1032));
  AND4_X1   g0832(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n959), .B2(new_n940), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1013), .A2(new_n1034), .ZN(G390));
  NAND4_X1  g0835(.A1(new_n731), .A2(G330), .A3(new_n815), .A4(new_n733), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n852), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n852), .B1(new_n886), .B2(new_n887), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1039), .A2(new_n895), .B1(new_n893), .B2(new_n891), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n812), .A2(new_n813), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n688), .B(new_n1041), .C1(new_n679), .C2(new_n715), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n811), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n852), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n878), .A3(new_n895), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT114), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n878), .A3(new_n1047), .A4(new_n895), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1038), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n891), .A2(new_n893), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT103), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n496), .B1(new_n655), .B2(new_n650), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n644), .B1(new_n1053), .B2(new_n703), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n663), .B(new_n667), .C1(new_n714), .C2(KEYINPUT26), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n687), .B(new_n814), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1052), .B1(new_n1056), .B2(new_n810), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n885), .A2(KEYINPUT103), .A3(new_n811), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1037), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1051), .B1(new_n1059), .B2(new_n896), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1038), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT115), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n882), .A2(new_n1063), .A3(G330), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1063), .B1(new_n882), .B2(G330), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n900), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1036), .B(new_n1037), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT116), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1069), .A2(new_n1043), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT116), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1068), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1050), .A2(new_n1062), .A3(new_n1067), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1067), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT117), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n707), .B(new_n1076), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n940), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1051), .A2(new_n792), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n244), .B1(new_n773), .B2(new_n312), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n825), .B1(new_n440), .B2(new_n749), .C1(new_n787), .C2(new_n745), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G107), .C2(new_n760), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n752), .A2(new_n214), .B1(new_n770), .B2(new_n371), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT118), .Z(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n784), .C2(new_n763), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT54), .B(G143), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(G125), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1091), .A2(new_n749), .B1(new_n1092), .B2(new_n763), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G128), .B2(new_n746), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n826), .B2(new_n752), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n244), .B(new_n1095), .C1(G159), .C2(new_n828), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n760), .A2(G137), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n218), .C2(new_n768), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n833), .A2(G150), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1089), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1101), .A2(new_n790), .B1(new_n279), .B2(new_n842), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1083), .A2(new_n741), .A3(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1082), .A2(KEYINPUT119), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT119), .B1(new_n1082), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1081), .B1(new_n1104), .B2(new_n1105), .ZN(G378));
  NAND2_X1  g0906(.A1(new_n1076), .A2(new_n1067), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT57), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n853), .B1(new_n890), .B2(new_n874), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n879), .C1(new_n1109), .C2(KEYINPUT40), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n433), .A2(new_n362), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT55), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n361), .A2(new_n858), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT56), .Z(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1112), .B(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1110), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n873), .A2(G330), .A3(new_n879), .A4(new_n1116), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n899), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n888), .A2(new_n897), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1122), .A2(new_n1118), .A3(new_n1119), .A4(new_n898), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1108), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1107), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n707), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT121), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT121), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1128), .A3(new_n707), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT122), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1076), .A2(new_n1067), .B1(new_n1123), .B2(new_n1121), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1107), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(KEYINPUT122), .A3(new_n1108), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1127), .A2(new_n1129), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n841), .A2(new_n218), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n759), .A2(new_n826), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G125), .A2(new_n746), .B1(new_n750), .B2(G137), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n355), .B2(new_n770), .C1(new_n773), .C2(new_n1091), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G128), .C2(new_n777), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT59), .ZN(new_n1142));
  AOI21_X1  g0942(.A(G41), .B1(new_n913), .B2(G124), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G33), .B1(new_n824), .B2(G159), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n218), .B1(new_n242), .B2(G41), .ZN(new_n1146));
  INV_X1    g0946(.A(G41), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n988), .A2(new_n1147), .A3(new_n244), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n770), .A2(new_n220), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n768), .A2(new_n276), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n745), .A2(new_n214), .B1(new_n763), .B2(new_n787), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(KEYINPUT120), .B1(new_n752), .B2(new_n445), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n752), .A2(KEYINPUT120), .A3(new_n445), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1153), .A2(new_n1154), .B1(new_n525), .B2(new_n750), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1152), .B(new_n1155), .C1(new_n440), .C2(new_n759), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT58), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1145), .A2(new_n1146), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n742), .B1(new_n1158), .B2(new_n790), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1137), .B(new_n1159), .C1(new_n1116), .C2(new_n793), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1133), .B2(new_n940), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1136), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G375));
  INV_X1    g0964(.A(new_n962), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1071), .A2(new_n1066), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  OR3_X1    g0967(.A1(new_n1079), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT123), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n1075), .A2(new_n940), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT124), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n745), .A2(new_n784), .B1(new_n752), .B2(new_n787), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n244), .B1(new_n763), .B2(new_n606), .C1(new_n371), .C2(new_n768), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G97), .C2(new_n833), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n750), .A2(G107), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n760), .A2(G116), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n990), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G159), .A2(new_n833), .B1(new_n913), .B2(G128), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT125), .Z(new_n1180));
  NAND2_X1  g0980(.A1(new_n760), .A2(new_n1090), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n770), .A2(new_n218), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n745), .A2(new_n826), .B1(new_n749), .B2(new_n355), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(G137), .C2(new_n777), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n307), .A3(new_n1181), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1178), .B1(new_n1185), .B2(new_n1150), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1186), .A2(new_n790), .B1(new_n220), .B2(new_n842), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n741), .B(new_n1187), .C1(new_n852), .C2(new_n793), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1075), .A2(KEYINPUT124), .A3(new_n940), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1172), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1169), .A2(new_n1191), .ZN(G381));
  NAND2_X1  g0992(.A1(new_n1082), .A2(new_n1103), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1081), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1163), .A2(new_n1196), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(G381), .A2(new_n1197), .A3(G384), .ZN(new_n1198));
  INV_X1    g0998(.A(G390), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n976), .A2(new_n978), .A3(new_n1199), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1200), .A2(G396), .A3(G393), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1201), .ZN(G407));
  OAI211_X1 g1002(.A(G407), .B(G213), .C1(G343), .C2(new_n1197), .ZN(G409));
  INV_X1    g1003(.A(KEYINPUT62), .ZN(new_n1204));
  INV_X1    g1004(.A(G213), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G343), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1075), .A2(new_n1067), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT60), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1166), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n708), .B1(new_n1166), .B2(new_n1208), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT126), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1213), .A2(KEYINPUT60), .A3(new_n1066), .A4(new_n1072), .ZN(new_n1214));
  AND4_X1   g1014(.A1(KEYINPUT126), .A2(new_n1214), .A3(new_n1211), .A4(new_n1077), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1191), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n845), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT126), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1077), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1211), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1210), .A2(KEYINPUT126), .A3(new_n1211), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G384), .A3(new_n1191), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1217), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1136), .A2(G378), .A3(new_n1162), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1162), .B1(new_n1134), .B2(new_n1165), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1196), .A2(new_n1227), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1206), .B(new_n1225), .C1(new_n1226), .C2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1204), .B1(new_n1229), .B2(KEYINPUT127), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1206), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G2897), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1217), .B(new_n1224), .C1(new_n1234), .C2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G384), .B1(new_n1223), .B2(new_n1191), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1190), .B(new_n845), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT61), .B1(new_n1233), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1225), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1231), .A2(new_n1232), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(KEYINPUT62), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1230), .A2(new_n1242), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n808), .B1(new_n983), .B2(new_n1010), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n975), .B2(G390), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n975), .A2(G390), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n975), .A2(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1200), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1250), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1253), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1247), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1253), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1240), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1244), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1229), .A2(KEYINPUT63), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1261), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1258), .A2(new_n1267), .ZN(G405));
  OAI21_X1  g1068(.A(new_n1226), .B1(new_n1163), .B2(new_n1195), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1243), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(new_n1243), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1257), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1257), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(G402));
endmodule


