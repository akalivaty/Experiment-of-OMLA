

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788;

  INV_X1 U370 ( .A(G953), .ZN(n779) );
  NOR2_X1 U371 ( .A1(n787), .A2(n788), .ZN(n424) );
  NAND2_X1 U372 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U373 ( .A(n764), .B(KEYINPUT71), .ZN(n525) );
  XNOR2_X1 U374 ( .A(n518), .B(n449), .ZN(n580) );
  XNOR2_X1 U375 ( .A(n560), .B(n350), .ZN(n537) );
  XOR2_X1 U376 ( .A(n524), .B(n523), .Z(n349) );
  XOR2_X1 U377 ( .A(KEYINPUT67), .B(KEYINPUT1), .Z(n350) );
  XNOR2_X2 U378 ( .A(n548), .B(n547), .ZN(n733) );
  XNOR2_X2 U379 ( .A(KEYINPUT92), .B(KEYINPUT18), .ZN(n454) );
  XNOR2_X2 U380 ( .A(G143), .B(G128), .ZN(n484) );
  BUF_X2 U381 ( .A(n742), .Z(n351) );
  XNOR2_X1 U382 ( .A(n535), .B(G472), .ZN(n742) );
  XNOR2_X2 U383 ( .A(n379), .B(G469), .ZN(n560) );
  INV_X1 U384 ( .A(n537), .ZN(n364) );
  NOR2_X1 U385 ( .A1(G953), .A2(G237), .ZN(n500) );
  XNOR2_X1 U386 ( .A(n777), .B(n522), .ZN(n533) );
  XNOR2_X1 U387 ( .A(n520), .B(n519), .ZN(n777) );
  XNOR2_X1 U388 ( .A(G128), .B(G110), .ZN(n511) );
  XNOR2_X1 U389 ( .A(n392), .B(G134), .ZN(n520) );
  INV_X1 U390 ( .A(KEYINPUT84), .ZN(n359) );
  NAND2_X1 U391 ( .A1(n443), .A2(n442), .ZN(n439) );
  AND2_X2 U392 ( .A1(n405), .A2(n572), .ZN(n404) );
  NOR2_X1 U393 ( .A1(n613), .A2(n426), .ZN(n425) );
  NAND2_X1 U394 ( .A1(n362), .A2(n361), .ZN(n360) );
  XNOR2_X1 U395 ( .A(n424), .B(KEYINPUT46), .ZN(n423) );
  XNOR2_X1 U396 ( .A(n623), .B(n622), .ZN(n787) );
  NAND2_X1 U397 ( .A1(n372), .A2(n373), .ZN(n709) );
  AND2_X1 U398 ( .A1(n726), .A2(n630), .ZN(n631) );
  XNOR2_X1 U399 ( .A(KEYINPUT41), .B(n625), .ZN(n757) );
  NOR2_X1 U400 ( .A1(n619), .A2(n624), .ZN(n621) );
  NOR2_X1 U401 ( .A1(n626), .A2(n396), .ZN(n609) );
  AND2_X1 U402 ( .A1(n582), .A2(n736), .ZN(n452) );
  INV_X1 U403 ( .A(n580), .ZN(n738) );
  NOR2_X1 U404 ( .A1(n692), .A2(G902), .ZN(n379) );
  XNOR2_X1 U405 ( .A(n418), .B(n776), .ZN(n686) );
  XNOR2_X1 U406 ( .A(n365), .B(n533), .ZN(n692) );
  XNOR2_X1 U407 ( .A(n515), .B(n419), .ZN(n418) );
  XNOR2_X1 U408 ( .A(n525), .B(n349), .ZN(n365) );
  XNOR2_X1 U409 ( .A(n513), .B(n420), .ZN(n419) );
  XNOR2_X1 U410 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U411 ( .A(n492), .B(n491), .ZN(n516) );
  XNOR2_X1 U412 ( .A(n456), .B(G146), .ZN(n492) );
  INV_X1 U413 ( .A(G953), .ZN(n389) );
  XNOR2_X1 U414 ( .A(G122), .B(KEYINPUT100), .ZN(n479) );
  XNOR2_X1 U415 ( .A(G143), .B(G128), .ZN(n392) );
  XOR2_X1 U416 ( .A(G110), .B(G104), .Z(n460) );
  XNOR2_X1 U417 ( .A(G101), .B(KEYINPUT68), .ZN(n390) );
  INV_X1 U418 ( .A(G125), .ZN(n456) );
  INV_X1 U419 ( .A(G953), .ZN(n388) );
  XNOR2_X1 U420 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  INV_X1 U421 ( .A(KEYINPUT88), .ZN(n363) );
  NAND2_X1 U422 ( .A1(n356), .A2(n352), .ZN(n362) );
  INV_X1 U423 ( .A(n353), .ZN(n352) );
  NAND2_X1 U424 ( .A1(n355), .A2(n354), .ZN(n353) );
  NAND2_X1 U425 ( .A1(n674), .A2(n359), .ZN(n354) );
  NAND2_X1 U426 ( .A1(n673), .A2(n359), .ZN(n355) );
  NAND2_X1 U427 ( .A1(n358), .A2(n357), .ZN(n356) );
  INV_X1 U428 ( .A(n674), .ZN(n357) );
  NOR2_X1 U429 ( .A1(n673), .A2(n359), .ZN(n358) );
  XNOR2_X2 U430 ( .A(n360), .B(KEYINPUT72), .ZN(n406) );
  AND2_X1 U431 ( .A1(n678), .A2(n554), .ZN(n361) );
  XNOR2_X1 U432 ( .A(n407), .B(n399), .ZN(n678) );
  XNOR2_X2 U433 ( .A(n546), .B(n545), .ZN(n674) );
  NOR2_X1 U434 ( .A1(n364), .A2(n736), .ZN(n737) );
  AND2_X1 U435 ( .A1(n558), .A2(n364), .ZN(n745) );
  NAND2_X1 U436 ( .A1(n452), .A2(n364), .ZN(n548) );
  XNOR2_X1 U437 ( .A(n537), .B(n363), .ZN(n587) );
  NOR2_X1 U438 ( .A1(n568), .A2(n364), .ZN(n569) );
  NAND2_X1 U439 ( .A1(n631), .A2(n537), .ZN(n633) );
  XNOR2_X2 U440 ( .A(n460), .B(G107), .ZN(n764) );
  XNOR2_X1 U441 ( .A(n367), .B(n366), .ZN(n459) );
  XNOR2_X1 U442 ( .A(n454), .B(n453), .ZN(n366) );
  XNOR2_X1 U443 ( .A(n484), .B(n521), .ZN(n367) );
  XNOR2_X1 U444 ( .A(n581), .B(KEYINPUT69), .ZN(n368) );
  NOR2_X2 U445 ( .A1(n637), .A2(n636), .ZN(n369) );
  NAND2_X1 U446 ( .A1(n609), .A2(KEYINPUT80), .ZN(n372) );
  NAND2_X1 U447 ( .A1(n370), .A2(n371), .ZN(n373) );
  INV_X1 U448 ( .A(n609), .ZN(n370) );
  INV_X1 U449 ( .A(KEYINPUT80), .ZN(n371) );
  INV_X1 U450 ( .A(n738), .ZN(n374) );
  XNOR2_X1 U451 ( .A(n581), .B(KEYINPUT69), .ZN(n604) );
  NOR2_X1 U452 ( .A1(n637), .A2(n636), .ZN(n778) );
  XNOR2_X2 U453 ( .A(n422), .B(KEYINPUT48), .ZN(n637) );
  XNOR2_X1 U454 ( .A(n469), .B(n398), .ZN(n375) );
  XNOR2_X1 U455 ( .A(n469), .B(n398), .ZN(n595) );
  INV_X1 U456 ( .A(n678), .ZN(n376) );
  INV_X1 U457 ( .A(n376), .ZN(n377) );
  INV_X1 U458 ( .A(n542), .ZN(n378) );
  XNOR2_X1 U459 ( .A(n351), .B(n541), .ZN(n582) );
  NAND2_X1 U460 ( .A1(n567), .A2(n380), .ZN(n539) );
  AND2_X1 U461 ( .A1(n374), .A2(n538), .ZN(n380) );
  NAND2_X1 U462 ( .A1(n769), .A2(n384), .ZN(n381) );
  NAND2_X1 U463 ( .A1(n381), .A2(n382), .ZN(n442) );
  OR2_X1 U464 ( .A1(n383), .A2(n448), .ZN(n382) );
  INV_X1 U465 ( .A(n402), .ZN(n383) );
  AND2_X1 U466 ( .A1(n778), .A2(n402), .ZN(n384) );
  NAND2_X1 U467 ( .A1(n567), .A2(n385), .ZN(n546) );
  AND2_X1 U468 ( .A1(n580), .A2(n543), .ZN(n385) );
  NAND2_X1 U469 ( .A1(n440), .A2(n439), .ZN(n386) );
  NAND2_X1 U470 ( .A1(n440), .A2(n439), .ZN(n438) );
  XNOR2_X2 U471 ( .A(n539), .B(KEYINPUT105), .ZN(n673) );
  NAND2_X1 U472 ( .A1(n406), .A2(n404), .ZN(n387) );
  NAND2_X1 U473 ( .A1(n406), .A2(n404), .ZN(n403) );
  XNOR2_X2 U474 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n453) );
  NAND2_X1 U475 ( .A1(n386), .A2(n644), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n387), .B(KEYINPUT45), .ZN(n393) );
  XNOR2_X1 U477 ( .A(n403), .B(KEYINPUT45), .ZN(n769) );
  NAND2_X1 U478 ( .A1(n641), .A2(n448), .ZN(n447) );
  XNOR2_X1 U479 ( .A(G104), .B(G122), .ZN(n496) );
  NAND2_X1 U480 ( .A1(n557), .A2(KEYINPUT44), .ZN(n405) );
  NOR2_X1 U481 ( .A1(n428), .A2(n432), .ZN(n431) );
  NAND2_X1 U482 ( .A1(n560), .A2(n435), .ZN(n437) );
  NAND2_X1 U483 ( .A1(n436), .A2(n435), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n410), .B(n409), .ZN(n408) );
  INV_X1 U485 ( .A(KEYINPUT34), .ZN(n409) );
  NAND2_X1 U486 ( .A1(n733), .A2(n550), .ZN(n410) );
  XNOR2_X1 U487 ( .A(KEYINPUT16), .B(G122), .ZN(n466) );
  AND2_X1 U488 ( .A1(n617), .A2(n603), .ZN(n427) );
  NAND2_X1 U489 ( .A1(n413), .A2(n394), .ZN(n412) );
  INV_X1 U490 ( .A(n636), .ZN(n413) );
  INV_X1 U491 ( .A(G237), .ZN(n468) );
  NOR2_X1 U492 ( .A1(n589), .A2(n578), .ZN(n429) );
  XOR2_X1 U493 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n527) );
  INV_X1 U494 ( .A(KEYINPUT10), .ZN(n491) );
  XNOR2_X1 U495 ( .A(G107), .B(G116), .ZN(n482) );
  XNOR2_X1 U496 ( .A(G140), .B(G113), .ZN(n494) );
  XNOR2_X1 U497 ( .A(KEYINPUT4), .B(G131), .ZN(n519) );
  NAND2_X1 U498 ( .A1(G237), .A2(G234), .ZN(n471) );
  INV_X1 U499 ( .A(G902), .ZN(n534) );
  XNOR2_X1 U500 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n464) );
  XNOR2_X1 U501 ( .A(n421), .B(KEYINPUT23), .ZN(n420) );
  INV_X1 U502 ( .A(G119), .ZN(n421) );
  AND2_X1 U503 ( .A1(G234), .A2(n388), .ZN(n485) );
  XNOR2_X1 U504 ( .A(n516), .B(n524), .ZN(n776) );
  NAND2_X1 U505 ( .A1(n438), .A2(n644), .ZN(n646) );
  XNOR2_X1 U506 ( .A(G140), .B(G137), .ZN(n524) );
  XNOR2_X1 U507 ( .A(KEYINPUT30), .B(KEYINPUT109), .ZN(n591) );
  INV_X1 U508 ( .A(n560), .ZN(n606) );
  INV_X1 U509 ( .A(n428), .ZN(n736) );
  XOR2_X1 U510 ( .A(n655), .B(KEYINPUT121), .Z(n656) );
  XOR2_X1 U511 ( .A(n647), .B(KEYINPUT59), .Z(n648) );
  XNOR2_X1 U512 ( .A(n662), .B(n665), .ZN(n666) );
  XNOR2_X1 U513 ( .A(n651), .B(KEYINPUT90), .ZN(n695) );
  NAND2_X1 U514 ( .A1(n408), .A2(n397), .ZN(n407) );
  AND2_X1 U515 ( .A1(n640), .A2(n447), .ZN(n394) );
  XOR2_X1 U516 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n395) );
  XOR2_X1 U517 ( .A(n416), .B(n395), .Z(n396) );
  XOR2_X1 U518 ( .A(n596), .B(n552), .Z(n397) );
  AND2_X1 U519 ( .A1(n470), .A2(G210), .ZN(n398) );
  XNOR2_X1 U520 ( .A(n553), .B(KEYINPUT35), .ZN(n399) );
  INV_X1 U521 ( .A(KEYINPUT76), .ZN(n435) );
  INV_X1 U522 ( .A(KEYINPUT65), .ZN(n642) );
  INV_X1 U523 ( .A(KEYINPUT82), .ZN(n448) );
  AND2_X1 U524 ( .A1(n638), .A2(n642), .ZN(n400) );
  AND2_X1 U525 ( .A1(n444), .A2(n642), .ZN(n401) );
  AND2_X1 U526 ( .A1(n394), .A2(KEYINPUT65), .ZN(n402) );
  NAND2_X1 U527 ( .A1(n411), .A2(n769), .ZN(n445) );
  NOR2_X1 U528 ( .A1(n637), .A2(n412), .ZN(n411) );
  XNOR2_X1 U529 ( .A(n391), .B(n645), .ZN(n414) );
  XNOR2_X1 U530 ( .A(n646), .B(n645), .ZN(n415) );
  XNOR2_X1 U531 ( .A(n646), .B(n645), .ZN(n690) );
  BUF_X1 U532 ( .A(n585), .Z(n416) );
  NAND2_X1 U533 ( .A1(n595), .A2(n726), .ZN(n585) );
  XNOR2_X1 U534 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U535 ( .A(n585), .B(n395), .ZN(n608) );
  XNOR2_X2 U536 ( .A(n562), .B(KEYINPUT103), .ZN(n712) );
  XNOR2_X2 U537 ( .A(n417), .B(n510), .ZN(n567) );
  NAND2_X2 U538 ( .A1(n549), .A2(n509), .ZN(n417) );
  XNOR2_X2 U539 ( .A(n478), .B(n477), .ZN(n549) );
  NAND2_X1 U540 ( .A1(n445), .A2(n401), .ZN(n441) );
  NAND2_X1 U541 ( .A1(n425), .A2(n423), .ZN(n422) );
  NAND2_X1 U542 ( .A1(n718), .A2(n427), .ZN(n426) );
  NAND2_X1 U543 ( .A1(n738), .A2(n739), .ZN(n428) );
  NAND2_X1 U544 ( .A1(n738), .A2(n429), .ZN(n436) );
  NAND2_X1 U545 ( .A1(n606), .A2(n736), .ZN(n590) );
  NAND2_X1 U546 ( .A1(n433), .A2(n430), .ZN(n594) );
  NAND2_X1 U547 ( .A1(n431), .A2(n606), .ZN(n430) );
  OR2_X1 U548 ( .A1(n589), .A2(n435), .ZN(n432) );
  AND2_X1 U549 ( .A1(n437), .A2(n434), .ZN(n433) );
  AND2_X2 U550 ( .A1(n441), .A2(n446), .ZN(n440) );
  NAND2_X1 U551 ( .A1(n643), .A2(n638), .ZN(n443) );
  NAND2_X1 U552 ( .A1(n394), .A2(KEYINPUT82), .ZN(n444) );
  NAND2_X1 U553 ( .A1(n643), .A2(n400), .ZN(n446) );
  NAND2_X1 U554 ( .A1(n608), .A2(n450), .ZN(n478) );
  XOR2_X1 U555 ( .A(KEYINPUT25), .B(n451), .Z(n449) );
  XOR2_X1 U556 ( .A(n476), .B(KEYINPUT95), .Z(n450) );
  AND2_X1 U557 ( .A1(n517), .A2(G217), .ZN(n451) );
  XNOR2_X1 U558 ( .A(n592), .B(n591), .ZN(n593) );
  INV_X1 U559 ( .A(KEYINPUT40), .ZN(n622) );
  INV_X1 U560 ( .A(KEYINPUT122), .ZN(n659) );
  XNOR2_X2 U561 ( .A(G101), .B(KEYINPUT68), .ZN(n521) );
  NAND2_X1 U562 ( .A1(n779), .A2(G224), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n455), .B(KEYINPUT87), .ZN(n457) );
  XNOR2_X1 U564 ( .A(n492), .B(n457), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n459), .B(n458), .ZN(n461) );
  XNOR2_X1 U566 ( .A(n461), .B(n525), .ZN(n467) );
  XNOR2_X1 U567 ( .A(G119), .B(G116), .ZN(n463) );
  XNOR2_X1 U568 ( .A(G113), .B(KEYINPUT70), .ZN(n462) );
  XNOR2_X1 U569 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U570 ( .A(n465), .B(n464), .ZN(n530) );
  XNOR2_X1 U571 ( .A(n530), .B(n466), .ZN(n766) );
  XNOR2_X1 U572 ( .A(n467), .B(n766), .ZN(n661) );
  NAND2_X1 U573 ( .A1(n661), .A2(n641), .ZN(n469) );
  NAND2_X1 U574 ( .A1(n534), .A2(n468), .ZN(n470) );
  NAND2_X1 U575 ( .A1(n470), .A2(G214), .ZN(n726) );
  XNOR2_X1 U576 ( .A(n471), .B(KEYINPUT14), .ZN(n474) );
  NAND2_X1 U577 ( .A1(G952), .A2(n474), .ZN(n472) );
  XOR2_X1 U578 ( .A(KEYINPUT93), .B(n472), .Z(n755) );
  NOR2_X1 U579 ( .A1(G953), .A2(n755), .ZN(n577) );
  NOR2_X1 U580 ( .A1(G898), .A2(n779), .ZN(n473) );
  XOR2_X1 U581 ( .A(KEYINPUT94), .B(n473), .Z(n767) );
  NAND2_X1 U582 ( .A1(G902), .A2(n474), .ZN(n573) );
  NOR2_X1 U583 ( .A1(n767), .A2(n573), .ZN(n475) );
  OR2_X1 U584 ( .A1(n577), .A2(n475), .ZN(n476) );
  INV_X1 U585 ( .A(KEYINPUT0), .ZN(n477) );
  XOR2_X1 U586 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n480) );
  XNOR2_X1 U587 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U588 ( .A(n481), .B(KEYINPUT101), .Z(n483) );
  XNOR2_X1 U589 ( .A(n483), .B(n482), .ZN(n488) );
  XNOR2_X1 U590 ( .A(KEYINPUT8), .B(n485), .ZN(n514) );
  NAND2_X1 U591 ( .A1(n514), .A2(G217), .ZN(n486) );
  XNOR2_X1 U592 ( .A(n520), .B(n486), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n655) );
  NAND2_X1 U594 ( .A1(n655), .A2(n534), .ZN(n490) );
  XOR2_X1 U595 ( .A(KEYINPUT102), .B(G478), .Z(n489) );
  XNOR2_X1 U596 ( .A(n490), .B(n489), .ZN(n563) );
  INV_X1 U597 ( .A(n563), .ZN(n551) );
  XNOR2_X1 U598 ( .A(n516), .B(KEYINPUT98), .ZN(n493) );
  XNOR2_X1 U599 ( .A(n493), .B(KEYINPUT11), .ZN(n504) );
  XOR2_X1 U600 ( .A(G131), .B(G143), .Z(n495) );
  XNOR2_X1 U601 ( .A(n495), .B(n494), .ZN(n499) );
  XOR2_X1 U602 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n497) );
  XNOR2_X1 U603 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U604 ( .A(n499), .B(n498), .ZN(n502) );
  XOR2_X1 U605 ( .A(KEYINPUT75), .B(n500), .Z(n526) );
  AND2_X1 U606 ( .A1(n526), .A2(G214), .ZN(n501) );
  XNOR2_X1 U607 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n504), .B(n503), .ZN(n647) );
  NAND2_X1 U609 ( .A1(n647), .A2(n534), .ZN(n506) );
  XOR2_X1 U610 ( .A(KEYINPUT13), .B(G475), .Z(n505) );
  XNOR2_X1 U611 ( .A(n506), .B(n505), .ZN(n564) );
  OR2_X1 U612 ( .A1(n551), .A2(n564), .ZN(n729) );
  NAND2_X1 U613 ( .A1(n641), .A2(G234), .ZN(n507) );
  XNOR2_X1 U614 ( .A(n507), .B(KEYINPUT20), .ZN(n517) );
  AND2_X1 U615 ( .A1(n517), .A2(G221), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n508), .B(KEYINPUT21), .ZN(n739) );
  INV_X1 U617 ( .A(n739), .ZN(n578) );
  NOR2_X1 U618 ( .A1(n729), .A2(n578), .ZN(n509) );
  XNOR2_X1 U619 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n510) );
  XOR2_X1 U620 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n512) );
  AND2_X1 U621 ( .A1(n514), .A2(G221), .ZN(n515) );
  NAND2_X1 U622 ( .A1(n686), .A2(n534), .ZN(n518) );
  XNOR2_X1 U623 ( .A(n390), .B(G146), .ZN(n522) );
  NAND2_X1 U624 ( .A1(n389), .A2(G227), .ZN(n523) );
  NAND2_X1 U625 ( .A1(n526), .A2(G210), .ZN(n529) );
  XNOR2_X1 U626 ( .A(n527), .B(G137), .ZN(n528) );
  XNOR2_X1 U627 ( .A(n529), .B(n528), .ZN(n531) );
  XNOR2_X1 U628 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U629 ( .A(n533), .B(n532), .ZN(n680) );
  NAND2_X1 U630 ( .A1(n680), .A2(n534), .ZN(n535) );
  INV_X1 U631 ( .A(n351), .ZN(n536) );
  AND2_X1 U632 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U633 ( .A(KEYINPUT104), .ZN(n540) );
  XNOR2_X1 U634 ( .A(n540), .B(KEYINPUT6), .ZN(n541) );
  INV_X1 U635 ( .A(n582), .ZN(n542) );
  AND2_X1 U636 ( .A1(n587), .A2(n542), .ZN(n543) );
  INV_X1 U637 ( .A(KEYINPUT66), .ZN(n544) );
  XNOR2_X1 U638 ( .A(n544), .B(KEYINPUT32), .ZN(n545) );
  XNOR2_X1 U639 ( .A(KEYINPUT86), .B(KEYINPUT33), .ZN(n547) );
  BUF_X1 U640 ( .A(n549), .Z(n550) );
  NAND2_X1 U641 ( .A1(n551), .A2(n564), .ZN(n596) );
  INV_X1 U642 ( .A(KEYINPUT79), .ZN(n552) );
  INV_X1 U643 ( .A(KEYINPUT78), .ZN(n553) );
  INV_X1 U644 ( .A(KEYINPUT44), .ZN(n554) );
  OR2_X1 U645 ( .A1(n673), .A2(n674), .ZN(n555) );
  INV_X1 U646 ( .A(n555), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n556), .A2(n377), .ZN(n557) );
  AND2_X1 U648 ( .A1(n736), .A2(n351), .ZN(n558) );
  NAND2_X1 U649 ( .A1(n550), .A2(n745), .ZN(n559) );
  XNOR2_X1 U650 ( .A(n559), .B(KEYINPUT31), .ZN(n715) );
  NOR2_X1 U651 ( .A1(n590), .A2(n351), .ZN(n561) );
  AND2_X1 U652 ( .A1(n550), .A2(n561), .ZN(n701) );
  OR2_X1 U653 ( .A1(n715), .A2(n701), .ZN(n566) );
  NAND2_X1 U654 ( .A1(n563), .A2(n564), .ZN(n562) );
  OR2_X1 U655 ( .A1(n564), .A2(n563), .ZN(n565) );
  INV_X1 U656 ( .A(n565), .ZN(n714) );
  NOR2_X1 U657 ( .A1(n712), .A2(n714), .ZN(n724) );
  INV_X1 U658 ( .A(n724), .ZN(n610) );
  NAND2_X1 U659 ( .A1(n566), .A2(n610), .ZN(n571) );
  BUF_X1 U660 ( .A(n567), .Z(n570) );
  OR2_X1 U661 ( .A1(n378), .A2(n374), .ZN(n568) );
  NAND2_X1 U662 ( .A1(n570), .A2(n569), .ZN(n698) );
  AND2_X1 U663 ( .A1(n571), .A2(n698), .ZN(n572) );
  NOR2_X1 U664 ( .A1(G900), .A2(n573), .ZN(n574) );
  NAND2_X1 U665 ( .A1(G953), .A2(n574), .ZN(n575) );
  XOR2_X1 U666 ( .A(KEYINPUT106), .B(n575), .Z(n576) );
  NOR2_X1 U667 ( .A1(n577), .A2(n576), .ZN(n589) );
  NOR2_X1 U668 ( .A1(n589), .A2(n578), .ZN(n579) );
  AND2_X1 U669 ( .A1(n712), .A2(n378), .ZN(n583) );
  NAND2_X1 U670 ( .A1(n368), .A2(n583), .ZN(n584) );
  XOR2_X1 U671 ( .A(KEYINPUT107), .B(n584), .Z(n629) );
  NOR2_X1 U672 ( .A1(n629), .A2(n416), .ZN(n586) );
  XNOR2_X1 U673 ( .A(n586), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n718) );
  NAND2_X1 U675 ( .A1(n726), .A2(n351), .ZN(n592) );
  NAND2_X1 U676 ( .A1(n594), .A2(n593), .ZN(n619) );
  INV_X1 U677 ( .A(n619), .ZN(n598) );
  INV_X1 U678 ( .A(n375), .ZN(n634) );
  NOR2_X1 U679 ( .A1(n596), .A2(n634), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n598), .A2(n597), .ZN(n671) );
  INV_X1 U681 ( .A(KEYINPUT81), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n671), .A2(n614), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n724), .A2(KEYINPUT47), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n671), .A2(n599), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n600), .A2(KEYINPUT81), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n603) );
  AND2_X1 U687 ( .A1(n604), .A2(n351), .ZN(n605) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT28), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n626) );
  NAND2_X1 U690 ( .A1(n709), .A2(n610), .ZN(n611) );
  NOR2_X1 U691 ( .A1(KEYINPUT47), .A2(n611), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT74), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n724), .A2(n614), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n709), .A2(n615), .ZN(n616) );
  NAND2_X1 U695 ( .A1(KEYINPUT47), .A2(n616), .ZN(n617) );
  INV_X1 U696 ( .A(KEYINPUT38), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n634), .B(n618), .ZN(n624) );
  XNOR2_X1 U698 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n621), .B(n620), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n628), .A2(n712), .ZN(n623) );
  INV_X1 U701 ( .A(n624), .ZN(n727) );
  NAND2_X1 U702 ( .A1(n727), .A2(n726), .ZN(n723) );
  NOR2_X1 U703 ( .A1(n723), .A2(n729), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n757), .A2(n626), .ZN(n627) );
  XNOR2_X1 U705 ( .A(KEYINPUT42), .B(n627), .ZN(n788) );
  NAND2_X1 U706 ( .A1(n628), .A2(n714), .ZN(n720) );
  INV_X1 U707 ( .A(n629), .ZN(n630) );
  XNOR2_X1 U708 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n633), .B(n632), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n672) );
  NAND2_X1 U711 ( .A1(n720), .A2(n672), .ZN(n636) );
  AND2_X2 U712 ( .A1(n393), .A2(n369), .ZN(n643) );
  INV_X1 U713 ( .A(n641), .ZN(n639) );
  AND2_X1 U714 ( .A1(KEYINPUT82), .A2(n639), .ZN(n638) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n721) );
  OR2_X1 U716 ( .A1(n641), .A2(n721), .ZN(n640) );
  BUF_X1 U717 ( .A(n643), .Z(n722) );
  NAND2_X1 U718 ( .A1(n722), .A2(KEYINPUT2), .ZN(n644) );
  INV_X1 U719 ( .A(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n415), .A2(G475), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(n652) );
  INV_X1 U722 ( .A(G952), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n650), .A2(G953), .ZN(n651) );
  NAND2_X1 U724 ( .A1(n652), .A2(n695), .ZN(n654) );
  INV_X1 U725 ( .A(KEYINPUT60), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(G60) );
  NAND2_X1 U727 ( .A1(n690), .A2(G478), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n658), .A2(n695), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G63) );
  NAND2_X1 U731 ( .A1(n415), .A2(G210), .ZN(n667) );
  BUF_X1 U732 ( .A(n661), .Z(n662) );
  XOR2_X1 U733 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n664) );
  XNOR2_X1 U734 ( .A(KEYINPUT85), .B(KEYINPUT55), .ZN(n663) );
  XOR2_X1 U735 ( .A(n664), .B(n663), .Z(n665) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n668), .A2(n695), .ZN(n670) );
  INV_X1 U738 ( .A(KEYINPUT56), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n670), .B(n669), .ZN(G51) );
  XNOR2_X1 U740 ( .A(n671), .B(G143), .ZN(G45) );
  XNOR2_X1 U741 ( .A(n672), .B(G140), .ZN(G42) );
  XOR2_X1 U742 ( .A(G110), .B(n673), .Z(G12) );
  BUF_X1 U743 ( .A(n674), .Z(n675) );
  XOR2_X1 U744 ( .A(G119), .B(KEYINPUT126), .Z(n676) );
  XNOR2_X1 U745 ( .A(n675), .B(n676), .ZN(G21) );
  XOR2_X1 U746 ( .A(G122), .B(KEYINPUT125), .Z(n677) );
  XNOR2_X1 U747 ( .A(n377), .B(n677), .ZN(G24) );
  NAND2_X1 U748 ( .A1(n414), .A2(G472), .ZN(n682) );
  XNOR2_X1 U749 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U751 ( .A1(n683), .A2(n695), .ZN(n685) );
  XOR2_X1 U752 ( .A(KEYINPUT89), .B(KEYINPUT63), .Z(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(G57) );
  NAND2_X1 U754 ( .A1(n690), .A2(G217), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n688), .A2(n695), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n689), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U758 ( .A1(n414), .A2(G469), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U760 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(n697) );
  INV_X1 U762 ( .A(n695), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(G54) );
  XOR2_X1 U764 ( .A(G101), .B(n698), .Z(n699) );
  XNOR2_X1 U765 ( .A(n699), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U766 ( .A1(n701), .A2(n712), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(G104), .ZN(G6) );
  XOR2_X1 U768 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U769 ( .A1(n701), .A2(n714), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U771 ( .A(G107), .B(n704), .ZN(G9) );
  XOR2_X1 U772 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n706) );
  NAND2_X1 U773 ( .A1(n714), .A2(n709), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n706), .B(n705), .ZN(n708) );
  XOR2_X1 U775 ( .A(G128), .B(KEYINPUT112), .Z(n707) );
  XNOR2_X1 U776 ( .A(n708), .B(n707), .ZN(G30) );
  NAND2_X1 U777 ( .A1(n709), .A2(n712), .ZN(n710) );
  XNOR2_X1 U778 ( .A(n710), .B(KEYINPUT114), .ZN(n711) );
  XNOR2_X1 U779 ( .A(G146), .B(n711), .ZN(G48) );
  NAND2_X1 U780 ( .A1(n715), .A2(n712), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n713), .B(G113), .ZN(G15) );
  NAND2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U783 ( .A(n716), .B(G116), .ZN(G18) );
  XNOR2_X1 U784 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U786 ( .A(G125), .B(n719), .ZN(G27) );
  XNOR2_X1 U787 ( .A(G134), .B(n720), .ZN(G36) );
  XNOR2_X1 U788 ( .A(n722), .B(n721), .ZN(n761) );
  NOR2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U790 ( .A(KEYINPUT117), .B(n725), .Z(n732) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U792 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U793 ( .A(KEYINPUT116), .B(n730), .ZN(n731) );
  NOR2_X1 U794 ( .A1(n732), .A2(n731), .ZN(n734) );
  INV_X1 U795 ( .A(n733), .ZN(n756) );
  NOR2_X1 U796 ( .A1(n734), .A2(n756), .ZN(n735) );
  XNOR2_X1 U797 ( .A(n735), .B(KEYINPUT118), .ZN(n751) );
  XOR2_X1 U798 ( .A(KEYINPUT50), .B(n737), .Z(n744) );
  NOR2_X1 U799 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U800 ( .A(KEYINPUT49), .B(n740), .Z(n741) );
  NOR2_X1 U801 ( .A1(n351), .A2(n741), .ZN(n743) );
  NAND2_X1 U802 ( .A1(n744), .A2(n743), .ZN(n747) );
  INV_X1 U803 ( .A(n745), .ZN(n746) );
  NAND2_X1 U804 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U805 ( .A(KEYINPUT51), .B(n748), .ZN(n749) );
  NOR2_X1 U806 ( .A1(n757), .A2(n749), .ZN(n750) );
  NOR2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U808 ( .A(n752), .B(KEYINPUT119), .Z(n753) );
  XNOR2_X1 U809 ( .A(KEYINPUT52), .B(n753), .ZN(n754) );
  NOR2_X1 U810 ( .A1(n755), .A2(n754), .ZN(n759) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n760) );
  OR2_X1 U813 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n762), .A2(G953), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n763), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U816 ( .A(n764), .B(G101), .Z(n765) );
  XNOR2_X1 U817 ( .A(n766), .B(n765), .ZN(n768) );
  NAND2_X1 U818 ( .A1(n768), .A2(n767), .ZN(n775) );
  AND2_X1 U819 ( .A1(n393), .A2(n388), .ZN(n773) );
  NAND2_X1 U820 ( .A1(G953), .A2(G224), .ZN(n770) );
  XNOR2_X1 U821 ( .A(KEYINPUT61), .B(n770), .ZN(n771) );
  AND2_X1 U822 ( .A1(n771), .A2(G898), .ZN(n772) );
  NOR2_X1 U823 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U824 ( .A(n775), .B(n774), .ZN(G69) );
  XNOR2_X1 U825 ( .A(n777), .B(n776), .ZN(n781) );
  XNOR2_X1 U826 ( .A(n369), .B(n781), .ZN(n780) );
  NAND2_X1 U827 ( .A1(n780), .A2(n389), .ZN(n786) );
  XOR2_X1 U828 ( .A(G227), .B(n781), .Z(n782) );
  XNOR2_X1 U829 ( .A(n782), .B(KEYINPUT124), .ZN(n783) );
  NAND2_X1 U830 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U831 ( .A1(G953), .A2(n784), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n786), .A2(n785), .ZN(G72) );
  XOR2_X1 U833 ( .A(G131), .B(n787), .Z(G33) );
  XOR2_X1 U834 ( .A(G137), .B(n788), .Z(G39) );
endmodule

