//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n467), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT66), .Z(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n461), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n474), .B(new_n478), .C1(G124), .C2(new_n481), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n466), .B2(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n484), .B(new_n487), .C1(new_n467), .C2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n461), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n481), .A2(G126), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n489), .A2(KEYINPUT67), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT67), .B1(new_n489), .B2(new_n493), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(G164));
  AND2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n503), .A2(new_n504), .B1(new_n497), .B2(new_n498), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n506), .A2(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT68), .Z(new_n515));
  INV_X1    g090(.A(new_n505), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n497), .A2(new_n498), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n515), .A2(new_n524), .ZN(G168));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n500), .A2(new_n526), .B1(new_n527), .B2(new_n505), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n511), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(G171));
  NOR2_X1   g106(.A1(new_n504), .A2(new_n503), .ZN(new_n532));
  INV_X1    g107(.A(G56), .ZN(new_n533));
  INV_X1    g108(.A(G68), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n519), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI221_X1 g112(.A(KEYINPUT69), .B1(new_n534), .B2(new_n519), .C1(new_n532), .C2(new_n533), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G651), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT71), .B(G81), .Z(new_n542));
  AOI22_X1  g117(.A1(new_n516), .A2(new_n542), .B1(new_n520), .B2(G43), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n539), .A2(new_n540), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n532), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(G651), .A2(new_n555), .B1(new_n516), .B2(G91), .ZN(new_n556));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n516), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n520), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n507), .B2(new_n508), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(G73), .A3(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n499), .A2(G86), .A3(new_n509), .ZN(new_n575));
  OAI211_X1 g150(.A(G48), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G305));
  INV_X1    g152(.A(G47), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT74), .B(G85), .Z(new_n579));
  OAI22_X1  g154(.A1(new_n500), .A2(new_n578), .B1(new_n505), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n511), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n580), .B2(new_n582), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n511), .B1(new_n500), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT76), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n516), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  AND2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n587), .B1(new_n594), .B2(G868), .ZN(G321));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G299), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G297));
  XOR2_X1   g174(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n476), .A2(G135), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT78), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  INV_X1    g184(.A(G111), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G2105), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(G123), .B2(new_n481), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT79), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2096), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(G2096), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2427), .ZN(new_n626));
  INV_X1    g201(.A(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT81), .B(G2438), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n626), .B(G2430), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n629), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(new_n633), .A3(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n634), .B(new_n637), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n642), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n646), .A3(G14), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g223(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n649), .B2(new_n654), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(new_n666), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  AND4_X1   g252(.A1(new_n672), .A2(new_n674), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n674), .A2(new_n676), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n677), .B1(new_n679), .B2(new_n672), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n664), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n663), .A3(new_n684), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(G29), .A2(G35), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G162), .B2(G29), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G2090), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT89), .B(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G20), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT23), .Z(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G299), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1956), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT102), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n696), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G19), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n546), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1341), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  INV_X1    g284(.A(G34), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT24), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(KEYINPUT24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G160), .B2(new_n709), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT95), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n462), .A2(G127), .ZN(new_n717));
  AND2_X1   g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  OAI21_X1  g293(.A(G2105), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n722));
  NAND2_X1  g297(.A1(G103), .A2(G2104), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G2105), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n476), .A2(G139), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n720), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G29), .B2(G33), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT94), .B(G2072), .Z(new_n731));
  AOI22_X1  g306(.A1(new_n716), .A2(G2084), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NOR2_X1   g308(.A1(G168), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n733), .B2(G21), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  NOR2_X1   g314(.A1(G29), .A2(G32), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT26), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n741), .B(new_n743), .C1(G141), .C2(new_n476), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G129), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT96), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(KEYINPUT97), .B(new_n740), .C1(new_n748), .C2(G29), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(new_n709), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(KEYINPUT97), .B2(new_n750), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n732), .B1(new_n738), .B2(KEYINPUT100), .C1(new_n739), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n709), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n476), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n481), .A2(G128), .ZN(new_n756));
  OR2_X1    g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n709), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n763), .B1(new_n735), .B2(new_n736), .C1(new_n615), .C2(new_n709), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT31), .B(G11), .Z(new_n765));
  XOR2_X1   g340(.A(KEYINPUT99), .B(G28), .Z(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT30), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G171), .A2(new_n733), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G5), .B2(new_n733), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n765), .B(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n773), .B1(new_n772), .B2(new_n771), .C1(new_n730), .C2(new_n731), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n752), .A2(new_n764), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n751), .A2(new_n739), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n778));
  NOR2_X1   g353(.A1(G164), .A2(new_n709), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G27), .B2(new_n709), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(G2078), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(G2078), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n715), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n778), .A2(new_n782), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n733), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n594), .B2(new_n733), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1348), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(G1348), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(new_n791), .C1(new_n694), .C2(G2090), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n701), .B2(new_n702), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n708), .A2(new_n775), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G23), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G288), .B2(new_n733), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT91), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT91), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n704), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n704), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n800), .A2(new_n801), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n709), .A2(G25), .ZN(new_n815));
  NOR2_X1   g390(.A1(G95), .A2(G2105), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT88), .Z(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n476), .A2(G131), .B1(G119), .B2(new_n481), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n709), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G24), .B(G290), .S(new_n704), .Z(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(G1986), .Z(new_n826));
  NAND4_X1  g401(.A1(new_n813), .A2(new_n814), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n794), .B1(new_n828), .B2(new_n829), .ZN(G311));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  INV_X1    g406(.A(new_n794), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(G150));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n532), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G651), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(KEYINPUT104), .A3(G651), .ZN(new_n840));
  AOI22_X1  g415(.A1(G93), .A2(new_n516), .B1(new_n520), .B2(G55), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n546), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n544), .A2(new_n545), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n842), .B(KEYINPUT105), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n591), .A2(new_n593), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n601), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n850), .A2(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n850), .A2(new_n852), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(KEYINPUT39), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n846), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(new_n747), .B(new_n759), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n489), .A2(new_n493), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n728), .ZN(new_n872));
  INV_X1    g447(.A(new_n869), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n868), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n727), .B(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n476), .A2(G142), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n461), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n481), .B2(G130), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(new_n619), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n821), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT108), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n872), .A2(new_n876), .A3(new_n885), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n614), .B(G160), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(G162), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(G162), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(KEYINPUT110), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT110), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n887), .B(new_n888), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n887), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n877), .A2(new_n886), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n891), .B(new_n890), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT109), .B(G37), .Z(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n846), .A2(new_n597), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n594), .A2(G299), .ZN(new_n902));
  INV_X1    g477(.A(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n851), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n848), .B(new_n603), .ZN(new_n910));
  MUX2_X1   g485(.A(new_n909), .B(new_n905), .S(new_n910), .Z(new_n911));
  XNOR2_X1  g486(.A(G290), .B(G305), .ZN(new_n912));
  XNOR2_X1  g487(.A(G166), .B(G288), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n911), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n901), .B1(new_n916), .B2(new_n597), .ZN(G295));
  OAI21_X1  g492(.A(new_n901), .B1(new_n916), .B2(new_n597), .ZN(G331));
  XNOR2_X1  g493(.A(G171), .B(KEYINPUT112), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G168), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n848), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n919), .B(G286), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n847), .A3(new_n844), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n909), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n905), .A3(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(new_n914), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n908), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n905), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(KEYINPUT41), .B2(new_n905), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n923), .B2(new_n921), .ZN(new_n936));
  INV_X1    g511(.A(new_n926), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n914), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n898), .A4(new_n928), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n932), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n928), .A2(new_n898), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n924), .B(new_n934), .C1(KEYINPUT41), .C2(new_n905), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n927), .B1(new_n944), .B2(new_n926), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT113), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n938), .A2(new_n947), .A3(new_n898), .A4(new_n928), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(KEYINPUT43), .A3(new_n948), .ZN(new_n949));
  OR3_X1    g524(.A1(new_n930), .A2(KEYINPUT43), .A3(new_n931), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n942), .B1(new_n951), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g527(.A(G125), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n464), .B1(new_n475), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G2105), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(G40), .A3(new_n469), .A4(new_n468), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n489), .B2(new_n493), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT45), .ZN(new_n958));
  INV_X1    g533(.A(G1996), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT46), .ZN(new_n961));
  INV_X1    g536(.A(new_n958), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n759), .B(new_n762), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(new_n748), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n747), .B(new_n959), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(new_n823), .A3(new_n821), .A4(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n760), .A2(new_n762), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n962), .A2(G290), .A3(G1986), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT48), .Z(new_n974));
  XOR2_X1   g549(.A(new_n821), .B(new_n823), .Z(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n963), .A3(new_n969), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n958), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n967), .A2(new_n968), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n980), .B(new_n981), .C1(new_n494), .C2(new_n495), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n869), .A2(new_n981), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n956), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1956), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n990));
  INV_X1    g565(.A(G91), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n990), .A2(new_n511), .B1(new_n991), .B2(new_n505), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT120), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n558), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(KEYINPUT120), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n556), .A2(KEYINPUT57), .A3(new_n558), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n556), .A2(KEYINPUT121), .A3(new_n558), .A4(KEYINPUT57), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n956), .B1(KEYINPUT45), .B2(new_n957), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT56), .B(G2072), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT67), .ZN(new_n1005));
  INV_X1    g580(.A(new_n488), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n487), .B1(new_n462), .B2(new_n484), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n490), .A2(new_n492), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n462), .A2(G2105), .ZN(new_n1010));
  INV_X1    g585(.A(G126), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1005), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n489), .A2(KEYINPUT67), .A3(new_n493), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1003), .B(new_n1004), .C1(new_n1015), .C2(KEYINPUT45), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n988), .A2(new_n1002), .A3(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n996), .A2(new_n1001), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1016), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n987), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n981), .B1(new_n494), .B2(new_n495), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n981), .B(new_n984), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n957), .A2(KEYINPUT115), .A3(new_n984), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G40), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n465), .A2(new_n1029), .A3(new_n470), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1348), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n983), .A2(new_n956), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n762), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n851), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1017), .B1(new_n1021), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT58), .B(G1341), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT45), .B(new_n981), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1030), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1022), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1039), .B1(new_n1043), .B2(new_n959), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n544), .A2(KEYINPUT122), .A3(new_n545), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1003), .B1(new_n1015), .B2(KEYINPUT45), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n1047), .A2(G1996), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1045), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1033), .A2(KEYINPUT60), .A3(new_n851), .A4(new_n1035), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1033), .A2(KEYINPUT60), .A3(new_n1035), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n594), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT60), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1052), .B(new_n1053), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1020), .A2(new_n1058), .A3(new_n1017), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1020), .B2(new_n1017), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1037), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1047), .A2(new_n804), .ZN(new_n1063));
  INV_X1    g638(.A(G2090), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1023), .A2(new_n1028), .A3(new_n1064), .A4(new_n1030), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G166), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT55), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(G8), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1030), .B2(new_n957), .ZN(new_n1071));
  INV_X1    g646(.A(G288), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G1976), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n570), .A2(new_n572), .ZN(new_n1082));
  OAI21_X1  g657(.A(G61), .B1(new_n504), .B2(new_n503), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n511), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G86), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n576), .B1(new_n505), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(G1981), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1981), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n574), .A2(new_n575), .A3(new_n1088), .A4(new_n576), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1081), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g667(.A(KEYINPUT116), .B(KEYINPUT49), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1087), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1080), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1096), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(KEYINPUT117), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1079), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n982), .A2(new_n986), .A3(new_n1064), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1043), .B2(G1971), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1069), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT119), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1106), .B(new_n1069), .C1(new_n1102), .C2(G8), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1070), .B(new_n1100), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1023), .A2(new_n1028), .A3(new_n784), .A4(new_n1030), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT45), .B(new_n981), .C1(new_n494), .C2(new_n495), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n956), .B1(new_n983), .B2(new_n1042), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n736), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1113), .A3(G168), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  AND2_X1   g690(.A1(KEYINPUT123), .A2(G8), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(G8), .A3(G286), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1115), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1108), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT124), .B(G1961), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1031), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1047), .B2(G2078), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(G2078), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1110), .A2(new_n1111), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G171), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1111), .A2(new_n1040), .A3(new_n1128), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1125), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(G171), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1130), .A2(G171), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1133), .B2(G171), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1062), .A2(new_n1123), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1067), .B1(new_n1063), .B2(new_n1101), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1106), .B1(new_n1140), .B2(new_n1069), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1103), .A2(KEYINPUT119), .A3(new_n1104), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1100), .A2(new_n1070), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1067), .B(G286), .C1(new_n1109), .C2(new_n1113), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1066), .A2(G8), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1104), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1144), .A2(KEYINPUT63), .A3(new_n1145), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1079), .B(new_n1070), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1071), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n1076), .A3(new_n1072), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1089), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1154), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(KEYINPUT118), .A3(new_n1089), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1153), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1108), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1121), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1119), .A4(new_n1117), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1131), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1139), .A2(new_n1152), .A3(new_n1161), .A4(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(G290), .B(G1986), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n958), .B1(new_n976), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1169), .A2(KEYINPUT125), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT125), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n979), .B1(new_n1172), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g749(.A1(G227), .A2(new_n459), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1176), .B1(new_n687), .B2(new_n689), .ZN(new_n1177));
  AND3_X1   g751(.A1(new_n1177), .A2(KEYINPUT127), .A3(new_n647), .ZN(new_n1178));
  AOI21_X1  g752(.A(KEYINPUT127), .B1(new_n1177), .B2(new_n647), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n899), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g754(.A1(new_n932), .A2(new_n940), .ZN(new_n1181));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1181), .ZN(G308));
  OR2_X1    g756(.A1(new_n1180), .A2(new_n1181), .ZN(G225));
endmodule


