

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  NOR2_X1 U323 ( .A1(n414), .A2(n419), .ZN(n420) );
  XNOR2_X1 U324 ( .A(n458), .B(KEYINPUT26), .ZN(n565) );
  XNOR2_X1 U325 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U326 ( .A(n446), .B(n445), .Z(n546) );
  XOR2_X1 U327 ( .A(KEYINPUT84), .B(G190GAT), .Z(n291) );
  AND2_X1 U328 ( .A1(G231GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U329 ( .A(n303), .B(G183GAT), .Z(n293) );
  XOR2_X1 U330 ( .A(n384), .B(n301), .Z(n294) );
  XNOR2_X1 U331 ( .A(n377), .B(n292), .ZN(n379) );
  XNOR2_X1 U332 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U333 ( .A(n361), .B(KEYINPUT76), .ZN(n362) );
  INV_X1 U334 ( .A(KEYINPUT98), .ZN(n465) );
  INV_X1 U335 ( .A(G78GAT), .ZN(n385) );
  XNOR2_X1 U336 ( .A(n363), .B(n362), .ZN(n366) );
  XNOR2_X1 U337 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U338 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U339 ( .A(KEYINPUT37), .B(n489), .ZN(n518) );
  XNOR2_X1 U340 ( .A(n374), .B(n373), .ZN(n414) );
  XOR2_X1 U341 ( .A(n308), .B(n307), .Z(n309) );
  XNOR2_X1 U342 ( .A(KEYINPUT38), .B(n492), .ZN(n501) );
  NOR2_X1 U343 ( .A1(n531), .A2(n449), .ZN(n453) );
  XNOR2_X1 U344 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U345 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT82), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U347 ( .A(KEYINPUT81), .B(G120GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U349 ( .A(KEYINPUT0), .B(n297), .Z(n425) );
  XOR2_X1 U350 ( .A(KEYINPUT20), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(G176GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n308) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G127GAT), .Z(n384) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G99GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n291), .B(n300), .ZN(n301) );
  NAND2_X1 U356 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n294), .B(n302), .ZN(n303) );
  XOR2_X1 U358 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n305) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n339) );
  XNOR2_X1 U361 ( .A(n339), .B(KEYINPUT83), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n293), .B(n306), .ZN(n307) );
  XOR2_X2 U363 ( .A(n425), .B(n309), .Z(n531) );
  XOR2_X1 U364 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n311) );
  XNOR2_X1 U365 ( .A(G211GAT), .B(G204GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U367 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n313) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n360) );
  XOR2_X1 U369 ( .A(G22GAT), .B(G155GAT), .Z(n377) );
  XNOR2_X1 U370 ( .A(n360), .B(n377), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U372 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U373 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U375 ( .A(n318), .B(KEYINPUT23), .Z(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n320) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n329), .B(KEYINPUT89), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n328) );
  XOR2_X1 U381 ( .A(G78GAT), .B(G148GAT), .Z(n324) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n355) );
  XOR2_X1 U384 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n326) );
  XNOR2_X1 U385 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n432) );
  XOR2_X1 U387 ( .A(n355), .B(n432), .Z(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n469) );
  XOR2_X1 U389 ( .A(n329), .B(KEYINPUT95), .Z(n331) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n332), .B(KEYINPUT94), .Z(n334) );
  XOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .Z(n368) );
  XNOR2_X1 U394 ( .A(G92GAT), .B(n368), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G204GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n335), .B(G64GAT), .ZN(n346) );
  XOR2_X1 U398 ( .A(n336), .B(n346), .Z(n341) );
  XOR2_X1 U399 ( .A(KEYINPUT78), .B(G211GAT), .Z(n338) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(G183GAT), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n381) );
  XNOR2_X1 U402 ( .A(n339), .B(n381), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n522) );
  XOR2_X1 U404 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n343) );
  NAND2_X1 U405 ( .A1(G230GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U407 ( .A(n344), .B(KEYINPUT70), .Z(n348) );
  XNOR2_X1 U408 ( .A(G71GAT), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n345), .B(KEYINPUT13), .ZN(n378) );
  XNOR2_X1 U410 ( .A(n346), .B(n378), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U412 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n350) );
  XNOR2_X1 U413 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U415 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U416 ( .A(KEYINPUT72), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U417 ( .A(G99GAT), .B(G85GAT), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n355), .B(n364), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n571) );
  XOR2_X1 U421 ( .A(G29GAT), .B(G43GAT), .Z(n359) );
  XNOR2_X1 U422 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n400) );
  XNOR2_X1 U424 ( .A(n360), .B(n400), .ZN(n363) );
  AND2_X1 U425 ( .A1(G232GAT), .A2(G233GAT), .ZN(n361) );
  XOR2_X1 U426 ( .A(n364), .B(KEYINPUT11), .Z(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(n368), .B(n367), .Z(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n370) );
  XNOR2_X1 U430 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n369) );
  XOR2_X1 U431 ( .A(n370), .B(n369), .Z(n372) );
  XNOR2_X1 U432 ( .A(G134GAT), .B(G218GAT), .ZN(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT36), .B(n414), .Z(n579) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n376) );
  XNOR2_X1 U435 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n390) );
  XOR2_X1 U437 ( .A(n380), .B(KEYINPUT14), .Z(n383) );
  XNOR2_X1 U438 ( .A(n381), .B(KEYINPUT80), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n388) );
  XNOR2_X1 U440 ( .A(G1GAT), .B(n384), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n390), .B(n389), .ZN(n486) );
  NOR2_X1 U442 ( .A1(n579), .A2(n486), .ZN(n391) );
  XOR2_X1 U443 ( .A(KEYINPUT45), .B(n391), .Z(n392) );
  NOR2_X1 U444 ( .A1(n571), .A2(n392), .ZN(n394) );
  INV_X1 U445 ( .A(KEYINPUT120), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n413) );
  XOR2_X1 U447 ( .A(G15GAT), .B(G22GAT), .Z(n396) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(G141GAT), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U450 ( .A(n397), .B(G36GAT), .Z(n399) );
  XOR2_X1 U451 ( .A(G113GAT), .B(G1GAT), .Z(n438) );
  XNOR2_X1 U452 ( .A(n438), .B(G50GAT), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n404) );
  XOR2_X1 U454 ( .A(n400), .B(KEYINPUT67), .Z(n402) );
  NAND2_X1 U455 ( .A1(G229GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U457 ( .A(n404), .B(n403), .Z(n412) );
  XOR2_X1 U458 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n406) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(G8GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U461 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n408) );
  XNOR2_X1 U462 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U465 ( .A(n412), .B(n411), .Z(n549) );
  INV_X1 U466 ( .A(n549), .ZN(n568) );
  NOR2_X1 U467 ( .A1(n413), .A2(n568), .ZN(n422) );
  XNOR2_X1 U468 ( .A(KEYINPUT117), .B(n486), .ZN(n561) );
  XOR2_X1 U469 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n416) );
  XOR2_X1 U470 ( .A(n571), .B(KEYINPUT41), .Z(n552) );
  NAND2_X1 U471 ( .A1(n552), .A2(n568), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  NOR2_X1 U473 ( .A1(n561), .A2(n417), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n418), .B(KEYINPUT119), .ZN(n419) );
  XOR2_X1 U475 ( .A(KEYINPUT47), .B(n420), .Z(n421) );
  NOR2_X1 U476 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n423), .B(KEYINPUT48), .ZN(n545) );
  NOR2_X1 U478 ( .A1(n522), .A2(n545), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n424), .B(KEYINPUT54), .ZN(n447) );
  INV_X1 U480 ( .A(n425), .ZN(n446) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n427) );
  XNOR2_X1 U482 ( .A(G57GAT), .B(KEYINPUT93), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n429) );
  XNOR2_X1 U485 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n431), .B(n430), .Z(n444) );
  XOR2_X1 U488 ( .A(n432), .B(KEYINPUT6), .Z(n434) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n442) );
  XOR2_X1 U491 ( .A(G155GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U492 ( .A(G127GAT), .B(G148GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n437), .B(G85GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U499 ( .A1(n447), .A2(n546), .ZN(n566) );
  NOR2_X1 U500 ( .A1(n469), .A2(n566), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  NAND2_X1 U502 ( .A1(n453), .A2(n414), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n450) );
  XOR2_X1 U504 ( .A(n552), .B(KEYINPUT109), .Z(n536) );
  NAND2_X1 U505 ( .A1(n536), .A2(n453), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(G176GAT), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NOR2_X1 U509 ( .A1(n571), .A2(n549), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT75), .B(n457), .Z(n490) );
  NAND2_X1 U511 ( .A1(n469), .A2(n531), .ZN(n458) );
  XOR2_X1 U512 ( .A(n522), .B(KEYINPUT27), .Z(n470) );
  INV_X1 U513 ( .A(n470), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n565), .A2(n459), .ZN(n548) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT96), .B(n460), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n531), .A2(n522), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n469), .A2(n461), .ZN(n462) );
  XOR2_X1 U519 ( .A(n463), .B(n462), .Z(n464) );
  NOR2_X1 U520 ( .A1(n548), .A2(n464), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n467), .A2(n546), .ZN(n473) );
  XOR2_X1 U523 ( .A(KEYINPUT28), .B(KEYINPUT64), .Z(n468) );
  XNOR2_X1 U524 ( .A(n469), .B(n468), .ZN(n527) );
  NAND2_X1 U525 ( .A1(n470), .A2(n527), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n546), .A2(n471), .ZN(n533) );
  NAND2_X1 U527 ( .A1(n531), .A2(n533), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n487) );
  OR2_X1 U529 ( .A1(n486), .A2(n414), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n474), .Z(n475) );
  AND2_X1 U531 ( .A1(n487), .A2(n475), .ZN(n508) );
  NAND2_X1 U532 ( .A1(n490), .A2(n508), .ZN(n484) );
  NOR2_X1 U533 ( .A1(n546), .A2(n484), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n522), .A2(n484), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT100), .B(n479), .Z(n480) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n480), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n531), .A2(n484), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U543 ( .A(G15GAT), .B(n483), .Z(G1326GAT) );
  NOR2_X1 U544 ( .A1(n527), .A2(n484), .ZN(n485) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  INV_X1 U546 ( .A(n486), .ZN(n575) );
  NOR2_X1 U547 ( .A1(n579), .A2(n575), .ZN(n488) );
  NAND2_X1 U548 ( .A1(n488), .A2(n487), .ZN(n489) );
  NAND2_X1 U549 ( .A1(n490), .A2(n518), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(KEYINPUT102), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n546), .A2(n501), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U554 ( .A(n495), .B(G29GAT), .Z(G1328GAT) );
  NOR2_X1 U555 ( .A1(n522), .A2(n501), .ZN(n496) );
  XOR2_X1 U556 ( .A(KEYINPUT104), .B(n496), .Z(n497) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U558 ( .A1(n531), .A2(n501), .ZN(n499) );
  XNOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U562 ( .A1(n527), .A2(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT111), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n549), .A2(n536), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT110), .B(n507), .Z(n519) );
  NAND2_X1 U571 ( .A1(n508), .A2(n519), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n546), .A2(n514), .ZN(n509) );
  XOR2_X1 U573 ( .A(n510), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n514), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT112), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U577 ( .A1(n531), .A2(n514), .ZN(n513) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n513), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n527), .A2(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT114), .ZN(n526) );
  NOR2_X1 U585 ( .A1(n526), .A2(n546), .ZN(n521) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n525) );
  NOR2_X1 U590 ( .A1(n531), .A2(n526), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  XNOR2_X1 U592 ( .A(KEYINPUT116), .B(KEYINPUT44), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n545), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n549), .A2(n535), .ZN(n534) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  INV_X1 U601 ( .A(n535), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n542), .A2(n536), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n540) );
  NAND2_X1 U605 ( .A1(n542), .A2(n561), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n414), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n551) );
  NOR2_X1 U613 ( .A1(n549), .A2(n551), .ZN(n550) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  INV_X1 U615 ( .A(n551), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n558), .A2(n552), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT122), .ZN(n554) );
  XOR2_X1 U618 ( .A(n554), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n558), .A2(n575), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n414), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n453), .A2(n568), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n453), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n570) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(n567), .B(KEYINPUT124), .Z(n578) );
  INV_X1 U634 ( .A(n578), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n574), .A2(n568), .ZN(n569) );
  XOR2_X1 U636 ( .A(n570), .B(n569), .Z(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n574), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT126), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

