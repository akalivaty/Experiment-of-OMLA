//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT66), .B(G238), .Z(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT67), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n213), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n207), .A2(G33), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT70), .ZN(new_n250));
  INV_X1    g0050(.A(G58), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n251), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n248), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(new_n207), .A3(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n202), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n248), .B1(G1), .B2(new_n207), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n202), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n258), .B2(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT74), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n276), .B1(new_n277), .B2(new_n274), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n213), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G274), .B1(new_n281), .B2(new_n213), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G41), .A2(G45), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G1), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n206), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n206), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(G226), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n283), .A2(new_n296), .A3(G190), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n283), .A2(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT76), .B1(new_n298), .B2(G200), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT76), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n300), .B(new_n301), .C1(new_n283), .C2(new_n296), .ZN(new_n302));
  OAI211_X1 g0102(.A(KEYINPUT75), .B(new_n297), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n272), .A2(new_n273), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n303), .B1(new_n270), .B2(new_n271), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n273), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  INV_X1    g0113(.A(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G33), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n315), .A2(new_n317), .A3(G226), .A4(new_n275), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n282), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n287), .A2(new_n288), .ZN(new_n321));
  INV_X1    g0121(.A(G274), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n293), .B2(new_n294), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n321), .A2(new_n323), .B1(new_n295), .B2(G238), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(new_n327), .A3(new_n324), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n311), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n320), .A2(new_n327), .A3(new_n324), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n327), .B1(new_n320), .B2(new_n324), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n329), .A2(new_n330), .B1(new_n333), .B2(G179), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n329), .B2(new_n330), .ZN(new_n336));
  OAI211_X1 g0136(.A(KEYINPUT77), .B(KEYINPUT14), .C1(new_n333), .C2(new_n311), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n250), .A2(G77), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n219), .A2(G20), .ZN(new_n340));
  INV_X1    g0140(.A(new_n256), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n340), .C1(new_n202), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT11), .A3(new_n247), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n206), .A2(KEYINPUT12), .A3(G13), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n340), .A2(new_n344), .B1(KEYINPUT12), .B2(new_n261), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n263), .B2(KEYINPUT12), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT11), .B1(new_n342), .B2(new_n247), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n333), .A2(G190), .ZN(new_n355));
  OAI21_X1  g0155(.A(G200), .B1(new_n331), .B2(new_n332), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n298), .A2(new_n311), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n283), .A2(new_n361), .A3(new_n296), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n266), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n365));
  INV_X1    g0165(.A(G107), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n365), .B1(new_n366), .B2(new_n274), .C1(new_n278), .C2(new_n220), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n282), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n289), .B1(G244), .B2(new_n295), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n364), .B1(new_n370), .B2(new_n311), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(G179), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n261), .A2(new_n277), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n263), .B2(new_n277), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G20), .A2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT72), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n376), .B1(new_n341), .B2(new_n253), .C1(new_n378), .C2(new_n249), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n375), .B1(new_n379), .B2(new_n247), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n372), .B2(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n373), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n370), .A2(G200), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n380), .C1(new_n384), .C2(new_n370), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n310), .A2(new_n359), .A3(new_n363), .A4(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n254), .A2(new_n261), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n254), .B2(new_n263), .ZN(new_n389));
  AND2_X1   g0189(.A1(KEYINPUT65), .A2(G68), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT65), .A2(G68), .ZN(new_n391));
  OAI21_X1  g0191(.A(G58), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n207), .B1(new_n392), .B2(new_n216), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n341), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT78), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT78), .ZN(new_n397));
  INV_X1    g0197(.A(new_n395), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n201), .B1(new_n218), .B2(G58), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n207), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n315), .A2(new_n317), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n402), .B2(new_n207), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  AOI211_X1 g0204(.A(new_n404), .B(G20), .C1(new_n315), .C2(new_n317), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n248), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n404), .B1(new_n274), .B2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n402), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n219), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n393), .A2(new_n395), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n412), .B2(KEYINPUT79), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n389), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n315), .A2(new_n317), .A3(G226), .A4(G1698), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n315), .A2(new_n317), .A3(G223), .A4(new_n275), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n282), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n321), .A2(new_n323), .B1(new_n295), .B2(G232), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n301), .ZN(new_n426));
  AND2_X1   g0226(.A1(KEYINPUT82), .A2(G190), .ZN(new_n427));
  NOR2_X1   g0227(.A1(KEYINPUT82), .A2(G190), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n426), .B1(new_n430), .B2(new_n425), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n418), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n389), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n398), .B1(new_n399), .B2(new_n207), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n218), .B1(new_n403), .B2(new_n405), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT79), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT16), .B1(new_n438), .B2(new_n413), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n396), .A2(new_n400), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n247), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n431), .B(new_n434), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(KEYINPUT83), .A2(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n433), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n423), .A2(new_n424), .A3(G179), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n311), .B1(new_n423), .B2(new_n424), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n425), .A2(G169), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n423), .A2(new_n424), .A3(G179), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n447), .B1(new_n418), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n451), .A2(new_n454), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n434), .B1(new_n439), .B2(new_n442), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT81), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n456), .A2(KEYINPUT18), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT18), .B1(new_n456), .B2(new_n459), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n446), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n387), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n315), .A2(new_n317), .A3(G264), .A4(G1698), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n315), .A2(new_n317), .A3(G257), .A4(new_n275), .ZN(new_n466));
  INV_X1    g0266(.A(G303), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n274), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n291), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT85), .B1(new_n472), .B2(new_n284), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n323), .A2(new_n474), .A3(new_n475), .A4(new_n469), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n468), .A2(new_n282), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT92), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n293), .A2(new_n294), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G270), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n472), .A2(KEYINPUT92), .A3(G270), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT93), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n477), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n477), .B2(new_n484), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n430), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n477), .A2(new_n484), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT93), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G200), .A3(new_n486), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n207), .C1(G33), .C2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n247), .C1(new_n207), .C2(G116), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT20), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n261), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G116), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n314), .A2(G1), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n261), .A2(new_n247), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n489), .A2(new_n492), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n311), .B1(new_n498), .B2(new_n503), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n491), .A2(new_n486), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n477), .A2(new_n484), .A3(G179), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n504), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n491), .A2(KEYINPUT21), .A3(new_n507), .A4(new_n486), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n506), .A2(new_n510), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n315), .A2(new_n317), .A3(new_n207), .A4(G68), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT89), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT89), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n274), .A2(new_n518), .A3(new_n207), .A4(G68), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n207), .B1(new_n313), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT88), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G87), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n494), .A3(new_n366), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT88), .B(new_n207), .C1(new_n313), .C2(new_n521), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n521), .B1(new_n249), .B2(new_n494), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n520), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT90), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n248), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n520), .A2(KEYINPUT90), .A3(new_n528), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n378), .A2(new_n261), .ZN(new_n535));
  INV_X1    g0335(.A(new_n378), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n282), .A2(new_n539), .A3(new_n469), .ZN(new_n540));
  OR2_X1    g0340(.A1(G238), .A2(G1698), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G244), .B2(new_n275), .ZN(new_n542));
  INV_X1    g0342(.A(G116), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n542), .A2(new_n402), .B1(new_n314), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n540), .B1(new_n544), .B2(new_n282), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n323), .A2(new_n469), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n323), .A2(new_n548), .A3(new_n469), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n311), .ZN(new_n552));
  INV_X1    g0352(.A(new_n551), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n361), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n538), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT91), .B1(new_n551), .B2(new_n384), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT91), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n545), .A2(new_n550), .A3(new_n557), .A4(G190), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n532), .A2(new_n533), .B1(new_n261), .B2(new_n378), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n502), .A2(G87), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n499), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n366), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n502), .A2(G107), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n315), .A2(new_n317), .A3(new_n207), .A4(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(KEYINPUT94), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n274), .A2(new_n207), .A3(G87), .A4(new_n572), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n314), .A2(new_n543), .A3(G20), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n207), .B2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n366), .A2(KEYINPUT23), .A3(G20), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n570), .B1(new_n586), .B2(new_n247), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n315), .A2(new_n317), .A3(G257), .A4(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n315), .A2(new_n317), .A3(G250), .A4(new_n275), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n479), .B1(new_n591), .B2(KEYINPUT95), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT95), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n588), .A2(new_n589), .A3(new_n593), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n473), .A2(new_n476), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n282), .B1(new_n469), .B2(new_n475), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G264), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n592), .A2(new_n594), .B1(G264), .B2(new_n597), .ZN(new_n601));
  AOI21_X1  g0401(.A(G200), .B1(new_n601), .B2(new_n596), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n587), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n315), .A2(new_n317), .A3(G250), .A4(G1698), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n315), .A2(new_n317), .A3(G244), .A4(new_n275), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT4), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n493), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n282), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n473), .A2(new_n476), .B1(new_n597), .B2(G257), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(G200), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n609), .A2(new_n610), .A3(G190), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n494), .A2(new_n366), .A3(KEYINPUT6), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT6), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n366), .A2(KEYINPUT84), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G107), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n617), .A2(new_n619), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n617), .A2(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n624));
  OAI21_X1  g0424(.A(G20), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n256), .A2(G77), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n366), .B1(new_n410), .B2(new_n411), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n247), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n499), .A2(G97), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n502), .B2(G97), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n615), .A2(new_n616), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n585), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n584), .B1(new_n576), .B2(new_n581), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n247), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n570), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n599), .A2(new_n311), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n601), .A2(new_n361), .A3(new_n596), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n609), .A2(new_n610), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n361), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n629), .A2(new_n631), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n611), .A2(new_n311), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n603), .A2(new_n633), .A3(new_n641), .A4(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n464), .A2(new_n515), .A3(new_n564), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n363), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n452), .A2(new_n453), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n458), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n382), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n354), .B1(new_n357), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n433), .A2(new_n445), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n657), .B2(new_n310), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n603), .A2(new_n633), .A3(new_n646), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n534), .A2(new_n561), .A3(new_n562), .A4(new_n535), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n560), .A2(KEYINPUT96), .A3(new_n561), .A4(new_n562), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n559), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n510), .A2(new_n641), .A3(new_n513), .A4(new_n514), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n659), .A2(new_n664), .A3(new_n555), .A4(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(new_n646), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n664), .A2(new_n667), .A3(new_n555), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n555), .A2(new_n563), .A3(new_n668), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT26), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n666), .A2(new_n669), .A3(new_n555), .A4(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n658), .B1(new_n464), .B2(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  INV_X1    g0478(.A(G213), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G343), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT97), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n505), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n515), .B2(new_n683), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n603), .A2(new_n641), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n587), .B2(new_n682), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n641), .B2(new_n682), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n682), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n641), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n675), .A2(new_n682), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n688), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n210), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n526), .A2(G116), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n217), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n642), .A2(new_n553), .A3(new_n601), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(new_n511), .ZN(new_n706));
  AOI21_X1  g0506(.A(G179), .B1(new_n545), .B2(new_n550), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(new_n611), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n491), .A3(new_n486), .A4(new_n599), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n611), .A2(new_n551), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n512), .A3(KEYINPUT30), .A4(new_n601), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n706), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT98), .B(KEYINPUT31), .Z(new_n713));
  AND3_X1   g0513(.A1(new_n712), .A2(new_n692), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n712), .B2(new_n692), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n489), .A2(new_n492), .A3(new_n505), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n675), .A2(new_n717), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n633), .A2(new_n603), .A3(new_n646), .A4(new_n641), .ZN(new_n719));
  INV_X1    g0519(.A(new_n564), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(new_n682), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT99), .B1(new_n722), .B2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT99), .ZN(new_n724));
  INV_X1    g0524(.A(G330), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n724), .B(new_n725), .C1(new_n716), .C2(new_n721), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n672), .A2(new_n682), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n670), .A2(KEYINPUT26), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n666), .A2(new_n731), .A3(new_n555), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n664), .A2(new_n555), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n667), .B1(new_n733), .B2(new_n668), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT29), .B(new_n682), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n703), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n685), .A2(G330), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n260), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n206), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n698), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n686), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT101), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n685), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n207), .B1(KEYINPUT102), .B2(new_n311), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n311), .A2(KEYINPUT102), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n213), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n207), .A2(new_n361), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n301), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n761), .A2(new_n346), .B1(new_n764), .B2(new_n277), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n762), .A2(new_n429), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(G58), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n301), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G20), .A3(G190), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n274), .B1(new_n769), .B2(new_n525), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n207), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(G107), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n394), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n759), .A2(new_n429), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n207), .B1(new_n775), .B2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n779), .A2(G50), .B1(G97), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n767), .A2(new_n774), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n769), .A2(new_n467), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n402), .B1(new_n772), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n776), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n784), .B(new_n786), .C1(G329), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n766), .A2(G322), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n760), .A2(new_n790), .B1(new_n763), .B2(G311), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n779), .A2(G326), .B1(G294), .B2(new_n781), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n757), .B1(new_n783), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n697), .A2(new_n402), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G355), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n210), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n697), .A2(new_n274), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n217), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n291), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n241), .A2(new_n291), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n756), .A2(new_n751), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n746), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n753), .A2(new_n794), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n748), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND3_X1  g0609(.A1(new_n373), .A2(new_n381), .A3(new_n682), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n380), .A2(new_n682), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(new_n385), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n810), .B1(new_n654), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n728), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n692), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n672), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n746), .B1(new_n727), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n727), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n756), .A2(new_n749), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n745), .B(new_n698), .C1(new_n277), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G294), .A2(new_n766), .B1(new_n763), .B2(G116), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n785), .B2(new_n761), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n402), .B1(new_n769), .B2(new_n366), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n772), .A2(new_n525), .B1(new_n776), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n779), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n827), .A2(new_n467), .B1(new_n494), .B2(new_n780), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n780), .A2(new_n251), .ZN(new_n830));
  INV_X1    g0630(.A(new_n769), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G50), .B1(new_n787), .B2(G132), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n832), .B(new_n274), .C1(new_n346), .C2(new_n772), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G137), .A2(new_n779), .B1(new_n763), .B2(G159), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  INV_X1    g0635(.A(new_n766), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n837), .C2(new_n761), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n830), .B(new_n833), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n813), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n821), .B1(new_n757), .B2(new_n842), .C1(new_n843), .C2(new_n750), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n819), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n743), .A2(new_n206), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n352), .A2(new_n692), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n353), .A2(new_n357), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n352), .B(new_n692), .C1(new_n338), .C2(new_n358), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n515), .A2(new_n647), .A3(new_n564), .A4(new_n692), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n712), .A2(new_n692), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n713), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n851), .B(new_n843), .C1(new_n852), .C2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT16), .B1(new_n401), .B2(new_n406), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n434), .B1(new_n858), .B2(new_n442), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n680), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n462), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n458), .A2(new_n680), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n443), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT37), .B1(new_n457), .B2(new_n458), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n859), .A2(new_n650), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n860), .A3(new_n443), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n862), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n418), .A2(new_n455), .A3(new_n447), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT81), .B1(new_n457), .B2(new_n458), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n652), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT18), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n656), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(KEYINPUT38), .B(new_n871), .C1(new_n877), .C2(new_n860), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n857), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n871), .B1(new_n877), .B2(new_n860), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n856), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT104), .B1(new_n887), .B2(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n863), .B1(new_n653), .B2(new_n446), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n651), .A2(new_n863), .A3(new_n443), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n865), .A2(new_n866), .B1(new_n891), .B2(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n885), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n857), .A2(new_n894), .A3(KEYINPUT40), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n713), .B1(new_n712), .B2(new_n692), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(KEYINPUT31), .B2(new_n854), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n721), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n463), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n725), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n896), .B2(new_n900), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n463), .A2(new_n730), .A3(new_n735), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n658), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT103), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n353), .A2(new_n692), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n816), .A2(new_n810), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n851), .C1(new_n872), .C2(new_n879), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n653), .A2(new_n680), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n905), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n847), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n902), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n623), .A2(new_n624), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n918), .A2(KEYINPUT35), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(KEYINPUT35), .ZN(new_n920));
  NOR4_X1   g0720(.A1(new_n919), .A2(new_n920), .A3(new_n543), .A4(new_n215), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT36), .Z(new_n922));
  NAND3_X1  g0722(.A1(new_n800), .A2(G77), .A3(new_n392), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n202), .A2(G68), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n260), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n917), .A2(new_n922), .A3(new_n926), .ZN(G367));
  AOI21_X1  g0727(.A(new_n805), .B1(new_n237), .B2(new_n798), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n210), .B2(new_n378), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n746), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n831), .A2(G116), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT46), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n931), .A2(new_n932), .B1(G303), .B2(new_n766), .ZN(new_n933));
  INV_X1    g0733(.A(G294), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n933), .B1(new_n366), .B2(new_n780), .C1(new_n934), .C2(new_n761), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n779), .A2(G311), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(new_n931), .B2(new_n932), .C1(new_n785), .C2(new_n764), .ZN(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n402), .B1(new_n776), .B2(new_n938), .C1(new_n494), .C2(new_n772), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT108), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n779), .A2(G143), .B1(G68), .B2(new_n781), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n837), .B2(new_n836), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT109), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G50), .A2(new_n763), .B1(new_n760), .B2(G159), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n773), .A2(G77), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n831), .A2(G58), .B1(new_n787), .B2(G137), .ZN(new_n949));
  AND4_X1   g0749(.A1(new_n274), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n930), .B1(new_n954), .B2(new_n756), .ZN(new_n955));
  INV_X1    g0755(.A(new_n555), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n560), .A2(new_n562), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n692), .ZN(new_n958));
  MUX2_X1   g0758(.A(new_n956), .B(new_n733), .S(new_n958), .Z(new_n959));
  OAI21_X1  g0759(.A(new_n955), .B1(new_n752), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n694), .A2(new_n688), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n690), .B2(new_n694), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(new_n686), .Z(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n738), .B2(new_n739), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n633), .B(new_n646), .C1(new_n632), .C2(new_n682), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n646), .B2(new_n682), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n695), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n695), .A2(new_n966), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n691), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n964), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n740), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n698), .B(KEYINPUT41), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n745), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n966), .B(KEYINPUT106), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n691), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT105), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n646), .B1(new_n979), .B2(new_n641), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n682), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n966), .A2(new_n688), .A3(new_n694), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT42), .Z(new_n987));
  AOI22_X1  g0787(.A1(new_n985), .A2(new_n987), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n983), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n960), .B1(new_n978), .B2(new_n989), .ZN(G387));
  OR3_X1    g0790(.A1(new_n964), .A2(KEYINPUT112), .A3(new_n699), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT112), .B1(new_n964), .B2(new_n699), .ZN(new_n992));
  INV_X1    g0792(.A(new_n963), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n992), .C1(new_n740), .C2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n690), .A2(new_n752), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n234), .A2(G45), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n253), .A2(G50), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT50), .Z(new_n998));
  OAI211_X1 g0798(.A(new_n700), .B(new_n291), .C1(new_n346), .C2(new_n277), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n996), .B(new_n798), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n700), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n795), .A2(new_n1001), .B1(new_n366), .B2(new_n697), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(KEYINPUT111), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n804), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT111), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n746), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G322), .A2(new_n779), .B1(new_n760), .B2(G311), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n467), .B2(new_n764), .C1(new_n938), .C2(new_n836), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT48), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n831), .A2(G294), .B1(new_n781), .B2(G283), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n772), .A2(new_n543), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n274), .B(new_n1017), .C1(G326), .C2(new_n787), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G50), .A2(new_n766), .B1(new_n763), .B2(G68), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n394), .B2(new_n827), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n831), .A2(G77), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n837), .B2(new_n776), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n402), .B(new_n1023), .C1(G97), .C2(new_n773), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n536), .A2(new_n781), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n760), .A2(new_n254), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1019), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1006), .B1(new_n1028), .B2(new_n756), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n993), .A2(new_n745), .B1(new_n995), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n994), .A2(new_n1030), .ZN(G393));
  AOI21_X1  g0831(.A(new_n699), .B1(new_n964), .B2(new_n973), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n964), .B2(new_n973), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n973), .A2(new_n745), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n799), .A2(new_n244), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n804), .B1(new_n494), .B2(new_n210), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n746), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G311), .A2(new_n766), .B1(new_n779), .B2(G317), .ZN(new_n1038));
  XOR2_X1   g0838(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n761), .A2(new_n467), .B1(new_n764), .B2(new_n934), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G116), .B2(new_n781), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n274), .B1(new_n773), .B2(G107), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n831), .A2(G283), .B1(new_n787), .B2(G322), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G150), .A2(new_n779), .B1(new_n766), .B2(G159), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n761), .A2(new_n202), .B1(new_n764), .B2(new_n253), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G77), .B2(new_n781), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n402), .B1(new_n773), .B2(G87), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n831), .A2(new_n218), .B1(new_n787), .B2(G143), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1045), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1037), .B1(new_n1053), .B2(new_n756), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n979), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n752), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1033), .A2(new_n1034), .A3(new_n1056), .ZN(G390));
  AOI21_X1  g0857(.A(new_n725), .B1(new_n898), .B2(new_n721), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1058), .A2(new_n843), .A3(new_n851), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n911), .A2(new_n851), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n909), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n907), .A2(new_n908), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n894), .A2(new_n1061), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n682), .B(new_n843), .C1(new_n732), .C2(new_n734), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n810), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n851), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1059), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n907), .A2(new_n908), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1065), .A2(new_n851), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n1061), .A3(new_n894), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n843), .B(new_n851), .C1(new_n723), .C2(new_n726), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n851), .B1(new_n1058), .B2(new_n843), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1065), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1073), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n843), .B1(new_n723), .B2(new_n726), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n851), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1059), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n911), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n463), .A2(new_n1058), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n903), .A2(new_n1084), .A3(new_n658), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1075), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1067), .A2(new_n1074), .A3(new_n1083), .A4(new_n1086), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n698), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1068), .A2(new_n749), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n820), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n746), .B1(new_n1093), .B2(new_n254), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n761), .A2(new_n366), .B1(new_n764), .B2(new_n494), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G116), .B2(new_n766), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n772), .A2(new_n346), .B1(new_n776), .B2(new_n934), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n274), .B(new_n1097), .C1(G87), .C2(new_n831), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n779), .A2(G283), .B1(G77), .B2(new_n781), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n274), .B1(new_n772), .B2(new_n202), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT114), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n769), .A2(new_n837), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n763), .A2(new_n1106), .B1(G159), .B2(new_n781), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G128), .A2(new_n779), .B1(new_n760), .B2(G137), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n766), .A2(G132), .B1(G125), .B2(new_n787), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1100), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT115), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n757), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1094), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1091), .A2(new_n745), .B1(new_n1092), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1090), .A2(new_n1116), .ZN(G378));
  NAND2_X1  g0917(.A1(new_n270), .A2(new_n680), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n310), .B2(new_n363), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1118), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n649), .B(new_n1120), .C1(new_n306), .C2(new_n309), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n308), .B1(new_n307), .B2(new_n273), .ZN(new_n1125));
  AND4_X1   g0925(.A1(new_n308), .A2(new_n272), .A3(new_n273), .A4(new_n304), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n363), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1120), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n310), .A2(new_n363), .A3(new_n1118), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n878), .A2(new_n893), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n843), .A4(new_n851), .ZN(new_n1134));
  OAI21_X1  g0934(.A(G330), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n889), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1131), .C1(new_n883), .C2(new_n888), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n914), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n887), .A2(KEYINPUT104), .A3(KEYINPUT40), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1131), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n914), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n889), .A2(new_n1136), .A3(new_n1132), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1089), .A2(new_n1086), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(KEYINPUT57), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n698), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT57), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1131), .A2(new_n749), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n746), .B1(new_n1093), .B2(G50), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n772), .A2(new_n251), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n274), .A2(G41), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1022), .A2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G283), .C2(new_n787), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n494), .A2(new_n761), .B1(new_n836), .B2(new_n366), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n827), .A2(new_n543), .B1(new_n346), .B2(new_n780), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1158), .B(new_n1161), .C1(new_n378), .C2(new_n764), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1163), .A2(KEYINPUT58), .B1(new_n1156), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT116), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(new_n1166), .B1(KEYINPUT58), .B2(new_n1163), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n779), .A2(G125), .B1(G150), .B2(new_n781), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT117), .Z(new_n1169));
  AOI22_X1  g0969(.A1(G132), .A2(new_n760), .B1(new_n763), .B2(G137), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n836), .C1(new_n769), .C2(new_n1105), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT118), .B(G124), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n787), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT59), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1177), .B1(new_n394), .B2(new_n772), .C1(new_n1173), .C2(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1154), .B1(new_n1180), .B2(new_n756), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1153), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1147), .B2(new_n745), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1152), .A2(new_n1184), .ZN(G375));
  OAI211_X1 g0985(.A(new_n1078), .B(new_n1085), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1087), .A2(new_n977), .A3(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT119), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n1080), .A2(new_n749), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n746), .B1(new_n1093), .B2(G68), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n779), .A2(G132), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT121), .Z(new_n1192));
  OAI22_X1  g0992(.A1(new_n769), .A2(new_n394), .B1(new_n776), .B2(new_n1171), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(new_n402), .A3(new_n1155), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n766), .A2(G137), .B1(G50), .B2(new_n781), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G150), .A2(new_n763), .B1(new_n760), .B2(new_n1106), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1025), .B1(new_n785), .B2(new_n836), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT120), .Z(new_n1199));
  AOI22_X1  g0999(.A1(new_n831), .A2(G97), .B1(new_n787), .B2(G303), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1200), .A2(new_n402), .A3(new_n948), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G107), .A2(new_n763), .B1(new_n760), .B2(G116), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n934), .C2(new_n827), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1197), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1190), .B1(new_n1204), .B2(new_n756), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1083), .A2(new_n745), .B1(new_n1189), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1188), .A2(new_n1206), .ZN(G381));
  NOR2_X1   g1007(.A1(G393), .A2(G396), .ZN(new_n1208));
  INV_X1    g1008(.A(G387), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  INV_X1    g1011(.A(G378), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n845), .A3(new_n1212), .ZN(new_n1213));
  OR4_X1    g1013(.A1(G375), .A2(new_n1210), .A3(G381), .A4(new_n1213), .ZN(G407));
  NOR2_X1   g1014(.A1(new_n679), .A2(G343), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(G375), .A2(G378), .A3(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT122), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1019(.A(KEYINPUT126), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1215), .A2(G2897), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1186), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT124), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n712), .A2(new_n692), .A3(new_n713), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n854), .B2(KEYINPUT31), .ZN(new_n1228));
  OAI21_X1  g1028(.A(G330), .B1(new_n852), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n724), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n722), .A2(KEYINPUT99), .A3(G330), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n851), .B1(new_n1232), .B2(new_n843), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n911), .B1(new_n1233), .B2(new_n1059), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1085), .B1(new_n1234), .B2(new_n1078), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1226), .B(new_n1186), .C1(new_n1235), .C2(new_n1222), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n699), .B1(new_n1224), .B2(KEYINPUT60), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1225), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1238), .A2(G384), .A3(new_n1206), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G384), .B1(new_n1238), .B2(new_n1206), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1221), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1206), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n845), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(G384), .A3(new_n1206), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1221), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1137), .A2(new_n1138), .A3(new_n914), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1144), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1148), .B(new_n977), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1147), .A2(new_n745), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1182), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1212), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT123), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1184), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1256), .A3(new_n1212), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1247), .B1(new_n1258), .B2(new_n1216), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1220), .B1(new_n1259), .B2(KEYINPUT61), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1256), .B1(new_n1252), .B2(new_n1212), .ZN(new_n1262));
  AOI211_X1 g1062(.A(KEYINPUT123), .B(G378), .C1(new_n1184), .C2(new_n1250), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1215), .B1(new_n1264), .B2(new_n1255), .ZN(new_n1265));
  OAI211_X1 g1065(.A(KEYINPUT126), .B(new_n1261), .C1(new_n1265), .C2(new_n1247), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1258), .A2(new_n1216), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(new_n1270), .A3(new_n1267), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1260), .A2(new_n1266), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1209), .A2(G390), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(new_n1211), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n808), .B1(new_n994), .B2(new_n1030), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1208), .B2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1208), .A2(new_n1276), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1247), .B1(new_n1265), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1258), .A2(new_n1216), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT125), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1268), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1267), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1280), .A2(KEYINPUT61), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1281), .A2(new_n1291), .ZN(G405));
  NOR2_X1   g1092(.A1(new_n1267), .A2(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1277), .B(new_n1279), .C1(KEYINPUT127), .C2(new_n1267), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1212), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1255), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(KEYINPUT127), .B2(new_n1267), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1296), .B(new_n1299), .ZN(G402));
endmodule


