//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G116), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(KEYINPUT69), .A3(G119), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT2), .B(G113), .Z(new_n195));
  AND2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  OR2_X1    g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n201), .A2(KEYINPUT0), .A3(G128), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n203), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(G134), .B2(new_n217), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n214), .A2(KEYINPUT11), .A3(G137), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(new_n215), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n213), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n206), .C2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G128), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT68), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n208), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n205), .A3(new_n207), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n217), .B2(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT66), .B1(new_n214), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n217), .A3(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n214), .A2(KEYINPUT67), .A3(G137), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n233), .A2(new_n223), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n225), .A2(new_n242), .A3(KEYINPUT30), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n203), .A2(new_n211), .A3(new_n212), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n244), .A2(KEYINPUT65), .B1(new_n223), .B2(new_n221), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n203), .A2(new_n211), .A3(new_n246), .A4(new_n212), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n241), .A2(new_n223), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n245), .A2(new_n247), .B1(new_n233), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n199), .B(new_n243), .C1(new_n249), .C2(KEYINPUT30), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n225), .A2(new_n242), .A3(new_n198), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT31), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(KEYINPUT28), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n258), .A2(KEYINPUT28), .ZN(new_n262));
  OAI22_X1  g076(.A1(new_n261), .A2(new_n262), .B1(new_n198), .B2(new_n249), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n256), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n258), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n224), .A3(new_n247), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT30), .B1(new_n268), .B2(new_n242), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n225), .A2(new_n242), .A3(KEYINPUT30), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n266), .B1(new_n271), .B2(new_n199), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n257), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n250), .A2(new_n274), .A3(new_n257), .A4(new_n258), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n265), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(G472), .A2(G902), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n187), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n225), .A2(new_n242), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n199), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n261), .B2(new_n262), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n263), .B2(new_n256), .ZN(new_n293));
  INV_X1    g107(.A(new_n272), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n256), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G472), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n259), .A2(KEYINPUT31), .B1(new_n263), .B2(new_n256), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n281), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n191), .B2(G128), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n230), .A2(KEYINPUT73), .A3(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n191), .A2(G128), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT24), .B(G110), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n191), .B2(G128), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT23), .A3(new_n306), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT23), .B1(new_n230), .B2(G119), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT74), .B1(new_n230), .B2(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n316), .B2(G110), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n320), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G146), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT77), .A4(G146), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n204), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n317), .A2(new_n326), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n307), .A2(new_n308), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT75), .B1(new_n316), .B2(G110), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n333));
  INV_X1    g147(.A(G110), .ZN(new_n334));
  AOI211_X1 g148(.A(new_n333), .B(new_n334), .C1(new_n312), .C2(new_n315), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n322), .A2(new_n323), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n204), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n324), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(KEYINPUT76), .A3(new_n204), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n330), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT78), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n330), .B(new_n348), .C1(new_n336), .C2(new_n342), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n282), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n350), .A2(KEYINPUT25), .A3(new_n282), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n282), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n350), .A2(new_n351), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT79), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n358), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n354), .B2(new_n355), .ZN(new_n365));
  INV_X1    g179(.A(new_n362), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n230), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n232), .B1(new_n370), .B2(new_n201), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G104), .ZN(new_n373));
  AND2_X1   g187(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n374));
  NOR2_X1   g188(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(G104), .A3(new_n372), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n376), .A2(new_n377), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(new_n381), .A3(KEYINPUT82), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n380), .A2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n386), .A3(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n371), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n382), .A2(new_n387), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n233), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n224), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT12), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G140), .ZN(new_n394));
  INV_X1    g208(.A(G227), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G953), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n394), .B(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n390), .A2(new_n391), .A3(new_n399), .A4(new_n224), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n382), .A2(KEYINPUT10), .A3(new_n387), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT10), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n401), .A2(new_n233), .B1(new_n388), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n224), .ZN(new_n404));
  OR2_X1    g218(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n384), .B1(new_n378), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n379), .A2(new_n381), .ZN(new_n407));
  OAI21_X1  g221(.A(G101), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n382), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n410), .B(G101), .C1(new_n406), .C2(new_n407), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n213), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n403), .A2(new_n404), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n393), .A2(new_n398), .A3(new_n400), .A4(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n403), .A2(new_n404), .A3(new_n412), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n404), .B1(new_n403), .B2(new_n412), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n397), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n282), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n393), .A2(new_n413), .A3(new_n400), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n397), .ZN(new_n422));
  OR3_X1    g236(.A1(new_n415), .A2(new_n416), .A3(new_n397), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G469), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n419), .A2(new_n282), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  OAI21_X1  g242(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT80), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n188), .A2(G122), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT92), .B1(new_n433), .B2(KEYINPUT14), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n188), .A2(G122), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n433), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n438));
  OAI21_X1  g252(.A(G107), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n206), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n230), .A2(G143), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G134), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n441), .A3(new_n214), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n433), .A3(new_n372), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(KEYINPUT91), .A3(new_n444), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n439), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n435), .A2(new_n433), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G107), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n448), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT13), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n440), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n206), .A2(KEYINPUT13), .A3(G128), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n455), .A2(new_n456), .A3(new_n441), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n453), .B(new_n444), .C1(new_n457), .C2(new_n214), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n428), .A2(new_n357), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n450), .A2(new_n458), .A3(new_n460), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(KEYINPUT87), .A2(G143), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G214), .A3(new_n252), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT87), .B(G143), .Z(new_n471));
  INV_X1    g285(.A(G237), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n344), .A3(G214), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n470), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT18), .A3(G131), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT18), .A2(G131), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n470), .B(new_n477), .C1(new_n471), .C2(new_n474), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n328), .B(new_n204), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT87), .A2(G143), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n469), .A2(new_n481), .B1(new_n252), .B2(G214), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n473), .A2(new_n468), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n470), .B(new_n222), .C1(new_n471), .C2(new_n474), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(KEYINPUT17), .A3(G131), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n480), .B1(new_n489), .B2(new_n342), .ZN(new_n490));
  XNOR2_X1  g304(.A(G113), .B(G122), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n380), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n342), .A2(new_n487), .A3(new_n488), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n492), .A4(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n340), .A2(new_n341), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n487), .A2(new_n488), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n492), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT90), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n493), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G475), .B1(new_n502), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT20), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n326), .A2(new_n327), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n484), .A2(new_n485), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n328), .B2(KEYINPUT89), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT19), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT19), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n328), .B2(new_n507), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n505), .B(new_n506), .C1(G146), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n492), .B1(new_n513), .B2(new_n496), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n495), .B1(new_n490), .B2(new_n492), .ZN(new_n516));
  AND4_X1   g330(.A1(new_n495), .A2(new_n494), .A3(new_n492), .A4(new_n496), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n504), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n514), .B1(new_n501), .B2(new_n497), .ZN(new_n521));
  INV_X1    g335(.A(new_n519), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n521), .A2(KEYINPUT20), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n467), .B(new_n503), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G214), .B1(G237), .B2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(G234), .A2(G237), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(G952), .A3(new_n344), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT21), .B(G898), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(G902), .A3(G953), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n532));
  XNOR2_X1  g346(.A(G110), .B(G122), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n537), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT8), .A3(new_n535), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n191), .A2(G116), .ZN(new_n543));
  OAI21_X1  g357(.A(G113), .B1(new_n543), .B2(KEYINPUT5), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n194), .A2(new_n195), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n382), .A4(new_n387), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n382), .A2(new_n387), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n196), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n541), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n549), .A2(new_n196), .A3(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n411), .B1(new_n196), .B2(new_n197), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n555), .B2(new_n409), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n539), .A2(new_n535), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n244), .A2(G125), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n229), .A2(new_n320), .A3(new_n232), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT7), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n344), .A2(G224), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT7), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n563), .B(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(G902), .B1(new_n558), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n382), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n548), .B1(new_n569), .B2(new_n554), .ZN(new_n570));
  INV_X1    g384(.A(new_n557), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n548), .B(new_n557), .C1(new_n569), .C2(new_n554), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(KEYINPUT6), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n559), .A2(new_n560), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n564), .B(KEYINPUT85), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT6), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n578), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G210), .B1(G237), .B2(G902), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n568), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n568), .B2(new_n580), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n525), .B(new_n531), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n432), .A2(new_n524), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n302), .A2(new_n369), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND2_X1  g401(.A1(new_n300), .A2(new_n282), .ZN(new_n588));
  INV_X1    g402(.A(G472), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT93), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n300), .A2(new_n282), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n414), .B2(new_n417), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n425), .B1(new_n594), .B2(new_n419), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n430), .B1(new_n595), .B2(new_n424), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n591), .A2(new_n369), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT94), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n503), .B1(new_n520), .B2(new_n523), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n465), .A2(new_n282), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n464), .B2(new_n465), .ZN(new_n601));
  INV_X1    g415(.A(new_n463), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n460), .B1(new_n450), .B2(new_n458), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT33), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n462), .A2(new_n605), .A3(new_n463), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n606), .A3(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n601), .A2(new_n607), .A3(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n599), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n584), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND3_X1  g431(.A1(new_n518), .A2(new_n504), .A3(new_n519), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT20), .B1(new_n521), .B2(new_n522), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n467), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(new_n503), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n584), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(KEYINPUT96), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n622), .B2(new_n584), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n598), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n343), .B(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n365), .B1(new_n361), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n432), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n524), .A2(new_n584), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n591), .A2(new_n635), .A3(new_n636), .A4(new_n593), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  OAI21_X1  g453(.A(new_n527), .B1(new_n530), .B2(G900), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AND4_X1   g456(.A1(new_n621), .A2(new_n620), .A3(new_n503), .A4(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n525), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n568), .A2(new_n580), .ZN(new_n645));
  INV_X1    g459(.A(new_n581), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n568), .A2(new_n580), .A3(new_n581), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT98), .B1(new_n643), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n525), .B1(new_n582), .B2(new_n583), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n622), .A2(new_n651), .A3(new_n652), .A4(new_n641), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n302), .B(new_n635), .C1(new_n650), .C2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NOR2_X1   g469(.A1(new_n582), .A2(new_n583), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n467), .B1(new_n620), .B2(new_n503), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n633), .A2(new_n361), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n359), .A2(new_n661), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n658), .A2(new_n660), .A3(new_n644), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n272), .A2(new_n256), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n284), .A2(new_n256), .A3(new_n258), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n282), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n281), .A2(new_n301), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n641), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n596), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n663), .A2(new_n668), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NAND3_X1  g488(.A1(new_n599), .A2(new_n612), .A3(new_n642), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n302), .A2(new_n649), .A3(new_n635), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  OR2_X1    g492(.A1(new_n594), .A2(new_n419), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(new_n431), .A3(new_n420), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n302), .A2(new_n369), .A3(new_n614), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n628), .A2(new_n302), .A3(new_n369), .A4(new_n680), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  XNOR2_X1  g499(.A(new_n594), .B(G469), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n649), .A2(new_n686), .A3(new_n431), .A4(new_n531), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n524), .A3(new_n634), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n302), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NAND2_X1  g504(.A1(new_n588), .A2(G472), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n285), .A2(new_n256), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n260), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n275), .A2(new_n277), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n259), .A2(KEYINPUT31), .B1(new_n285), .B2(new_n256), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n279), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n365), .A2(new_n366), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n691), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n680), .A2(new_n659), .A3(new_n649), .A4(new_n531), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT101), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n687), .A2(new_n660), .ZN(new_n705));
  AOI22_X1  g519(.A1(G472), .A2(new_n588), .B1(new_n699), .B2(new_n279), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n707), .A4(new_n701), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  NAND2_X1  g524(.A1(new_n686), .A2(new_n431), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n651), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n706), .A2(new_n662), .A3(new_n676), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  NOR3_X1   g528(.A1(new_n582), .A2(new_n583), .A3(new_n644), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n596), .B2(KEYINPUT102), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n432), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT103), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n647), .A2(new_n525), .A3(new_n648), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n432), .B2(new_n717), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n596), .A2(KEYINPUT102), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n675), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n302), .A2(KEYINPUT104), .A3(new_n701), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT104), .B1(new_n302), .B2(new_n701), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n719), .A2(new_n724), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n359), .A2(KEYINPUT79), .A3(new_n362), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n367), .B1(new_n365), .B2(new_n366), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n187), .B(new_n280), .C1(new_n695), .C2(new_n297), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT32), .B1(new_n300), .B2(new_n279), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n732), .B1(new_n735), .B2(new_n296), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n728), .A2(KEYINPUT42), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n643), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n729), .A2(new_n736), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT106), .B(G134), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G36));
  AOI21_X1  g559(.A(new_n599), .B1(new_n610), .B2(new_n611), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT43), .ZN(new_n747));
  AOI211_X1 g561(.A(G902), .B(new_n590), .C1(new_n695), .C2(new_n297), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n592), .B1(new_n300), .B2(new_n282), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n751), .A3(new_n662), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n720), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n422), .A2(new_n423), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n419), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT107), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n425), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n420), .B1(new_n762), .B2(KEYINPUT46), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n431), .B(new_n669), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n756), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT108), .B(G137), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G39));
  OAI21_X1  g583(.A(new_n431), .B1(new_n763), .B2(new_n764), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT47), .B(new_n431), .C1(new_n763), .C2(new_n764), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n302), .A2(new_n369), .A3(new_n675), .A4(new_n720), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND2_X1  g591(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n737), .A2(new_n738), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n302), .A2(new_n369), .A3(new_n680), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n628), .A2(new_n781), .B1(new_n704), .B2(new_n708), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  INV_X1    g597(.A(new_n586), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n613), .A2(new_n622), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n624), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n637), .B1(new_n597), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n681), .A2(new_n689), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n584), .B1(new_n613), .B2(new_n622), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n596), .A2(new_n731), .A3(new_n730), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n750), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n586), .A2(new_n794), .A3(KEYINPUT111), .A4(new_n637), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n782), .A2(new_n788), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n780), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n697), .A2(new_n696), .B1(new_n275), .B2(new_n277), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n280), .B1(new_n798), .B2(new_n694), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n589), .B1(new_n300), .B2(new_n282), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n799), .A2(new_n675), .A3(new_n800), .A4(new_n634), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n729), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n662), .A2(new_n431), .A3(new_n427), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n735), .B2(new_n296), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n647), .A2(new_n525), .A3(new_n648), .A4(new_n642), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n524), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT112), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(KEYINPUT113), .A2(new_n743), .A3(new_n802), .A4(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n801), .A2(new_n729), .B1(new_n804), .B2(new_n807), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT113), .B1(new_n810), .B2(new_n743), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n659), .A2(new_n649), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n596), .A2(new_n634), .A3(new_n642), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n668), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n654), .A2(new_n677), .A3(new_n713), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT52), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n797), .A2(KEYINPUT53), .A3(new_n812), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n792), .A2(new_n748), .A3(new_n749), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n803), .A2(new_n524), .A3(new_n584), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n824), .A2(new_n791), .B1(new_n750), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT111), .B1(new_n826), .B2(new_n586), .ZN(new_n827));
  AND4_X1   g641(.A1(KEYINPUT111), .A2(new_n586), .A3(new_n637), .A4(new_n794), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n701), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n799), .A2(new_n800), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n707), .B1(new_n831), .B2(new_n705), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n702), .A2(KEYINPUT101), .A3(new_n703), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n684), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n789), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n739), .A2(new_n829), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n743), .A2(new_n802), .A3(new_n808), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n810), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n817), .B(KEYINPUT52), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n836), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n822), .B(new_n823), .C1(new_n843), .C2(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n836), .A2(new_n841), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n847), .B2(new_n821), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n844), .B1(new_n850), .B2(new_n823), .ZN(new_n851));
  INV_X1    g665(.A(G952), .ZN(new_n852));
  INV_X1    g666(.A(new_n527), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n747), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n831), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n852), .B(G953), .C1(new_n855), .C2(new_n712), .ZN(new_n856));
  INV_X1    g670(.A(new_n668), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n711), .A2(new_n720), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n369), .A3(new_n853), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n726), .A2(new_n727), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n862), .B2(new_n863), .ZN(new_n866));
  OAI221_X1 g680(.A(new_n856), .B1(new_n613), .B2(new_n859), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n855), .A2(new_n644), .A3(new_n658), .A4(new_n680), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT50), .Z(new_n869));
  AND2_X1   g683(.A1(new_n686), .A2(new_n430), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n715), .B(new_n855), .C1(new_n774), .C2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n854), .A2(new_n662), .A3(new_n706), .A4(new_n858), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n859), .A2(new_n599), .A3(new_n612), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n869), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n867), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n851), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n830), .A2(new_n430), .A3(new_n644), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n879), .B(new_n746), .C1(new_n880), .C2(new_n686), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT109), .Z(new_n882));
  INV_X1    g696(.A(new_n658), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n880), .B2(new_n686), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n857), .A3(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT110), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n878), .A2(new_n886), .ZN(G75));
  OAI21_X1  g701(.A(new_n822), .B1(new_n843), .B2(KEYINPUT53), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(G902), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n574), .A2(new_n579), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n577), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n852), .A2(G953), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT117), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n895), .A2(new_n896), .A3(new_n899), .ZN(G51));
  NAND2_X1  g714(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(KEYINPUT118), .A3(new_n844), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n888), .A2(new_n903), .A3(KEYINPUT54), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n425), .B(KEYINPUT57), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT119), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n902), .A2(new_n908), .A3(new_n904), .A4(new_n905), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n418), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n889), .A2(new_n761), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n899), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n521), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n898), .B1(new_n913), .B2(new_n521), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n913), .B2(new_n521), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n604), .A2(new_n606), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n600), .B(KEYINPUT59), .Z(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n851), .B2(new_n920), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n919), .A2(new_n902), .A3(new_n904), .A4(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n899), .A3(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  AND2_X1   g739(.A1(new_n888), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n633), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n927), .B(new_n898), .C1(new_n360), .C2(new_n926), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT61), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G66));
  INV_X1    g745(.A(G224), .ZN(new_n932));
  OAI21_X1  g746(.A(G953), .B1(new_n528), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n796), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n892), .B1(G898), .B2(new_n344), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT122), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  AOI22_X1  g752(.A1(new_n774), .A2(new_n775), .B1(new_n756), .B2(new_n766), .ZN(new_n939));
  INV_X1    g753(.A(new_n670), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n736), .A2(new_n940), .A3(new_n715), .A4(new_n785), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n654), .A2(new_n677), .A3(new_n713), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT123), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n673), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n943), .A3(new_n673), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT124), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n271), .B(new_n512), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n344), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n861), .A2(new_n813), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n766), .A2(new_n953), .B1(new_n737), .B2(new_n742), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n939), .A2(new_n945), .A3(new_n739), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n344), .ZN(new_n956));
  INV_X1    g770(.A(G900), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n951), .B1(new_n957), .B2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n395), .B2(new_n957), .ZN(new_n959));
  AOI22_X1  g773(.A1(new_n956), .A2(new_n958), .B1(KEYINPUT125), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n952), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G72));
  NOR2_X1   g777(.A1(new_n294), .A2(new_n257), .ZN(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n964), .A2(new_n664), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n955), .B2(new_n796), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n964), .B1(new_n969), .B2(KEYINPUT127), .ZN(new_n971));
  OAI221_X1 g785(.A(new_n898), .B1(new_n850), .B2(new_n968), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n947), .A2(new_n934), .A3(new_n949), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n664), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n973), .B2(new_n966), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n972), .A2(new_n978), .ZN(G57));
endmodule


