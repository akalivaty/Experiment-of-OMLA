//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n206));
  NAND2_X1  g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G218gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT72), .B1(new_n214), .B2(new_n207), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n208), .B2(new_n209), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(KEYINPUT72), .A3(new_n207), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT73), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT71), .A3(new_n220), .ZN(new_n224));
  OR2_X1    g023(.A1(G197gat), .A2(G204gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G197gat), .A2(G204gat), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n223), .A2(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n216), .A2(new_n219), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(new_n224), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT71), .B1(new_n207), .B2(new_n220), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n218), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n206), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238));
  NAND2_X1  g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239));
  INV_X1    g038(.A(G155gat), .ZN(new_n240));
  INV_X1    g039(.A(G162gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G141gat), .B(G148gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n239), .B(new_n242), .C1(new_n243), .C2(KEYINPUT2), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  INV_X1    g044(.A(G148gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT75), .B(G148gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n249), .B2(G141gat), .ZN(new_n250));
  OR2_X1    g049(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n251), .A2(KEYINPUT76), .A3(G141gat), .A4(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n239), .B1(new_n242), .B2(KEYINPUT2), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n238), .B(new_n244), .C1(new_n250), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n236), .B1(new_n237), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G141gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n248), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n253), .B(new_n254), .C1(new_n260), .C2(new_n247), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n244), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n228), .A2(new_n237), .A3(new_n234), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT3), .B1(new_n264), .B2(KEYINPUT81), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n228), .A2(new_n234), .A3(new_n266), .A4(new_n237), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n258), .B1(new_n268), .B2(KEYINPUT82), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT82), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n270), .B(new_n263), .C1(new_n265), .C2(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n205), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G22gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n236), .A2(new_n237), .A3(new_n262), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n238), .B1(new_n261), .B2(new_n244), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(new_n205), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(new_n272), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT83), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n264), .A2(KEYINPUT81), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n238), .A3(new_n267), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n262), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n257), .B1(new_n283), .B2(new_n270), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n204), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n277), .ZN(new_n287));
  OAI21_X1  g086(.A(G22gat), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G78gat), .B(G106gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT31), .B(G50gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT67), .A2(KEYINPUT34), .ZN(new_n297));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G113gat), .ZN(new_n300));
  INV_X1    g099(.A(G113gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n306));
  NOR2_X1   g105(.A1(G127gat), .A2(G134gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G127gat), .A2(G134gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n309), .ZN(new_n312));
  OAI22_X1  g111(.A1(new_n312), .A2(new_n307), .B1(KEYINPUT65), .B2(KEYINPUT1), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(new_n300), .B2(new_n302), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n319), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n318), .A2(G169gat), .A3(G176gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT64), .B1(new_n320), .B2(new_n323), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n324), .A2(KEYINPUT64), .A3(KEYINPUT25), .A4(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(G169gat), .ZN(new_n334));
  INV_X1    g133(.A(G176gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n322), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(KEYINPUT28), .A3(new_n340), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n317), .B1(new_n332), .B2(new_n346), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n316), .B(new_n345), .C1(new_n330), .C2(new_n331), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n298), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(KEYINPUT67), .A2(KEYINPUT34), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n297), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n347), .B2(new_n348), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT64), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n324), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n355), .A2(KEYINPUT25), .B1(new_n324), .B2(new_n326), .ZN(new_n356));
  INV_X1    g155(.A(new_n331), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n346), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n316), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n332), .A2(new_n317), .A3(new_n346), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT68), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n361), .A3(new_n298), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT66), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n359), .A2(G227gat), .A3(G233gat), .A4(new_n360), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(KEYINPUT32), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n364), .A3(KEYINPUT32), .ZN(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n365), .B(KEYINPUT32), .C1(new_n372), .C2(new_n371), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n363), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n368), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n375), .B(new_n363), .C1(new_n377), .C2(new_n366), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT69), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n374), .A2(new_n380), .A3(new_n375), .A4(new_n363), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n294), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n316), .A2(new_n261), .A3(new_n244), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n316), .A2(new_n261), .A3(KEYINPUT4), .A4(new_n244), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n311), .A2(KEYINPUT77), .A3(new_n315), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT77), .B1(new_n311), .B2(new_n315), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n256), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n386), .B(new_n387), .C1(new_n390), .C2(new_n275), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n392), .B(KEYINPUT78), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n262), .B1(new_n388), .B2(new_n389), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n384), .ZN(new_n396));
  OAI22_X1  g195(.A1(new_n391), .A2(new_n393), .B1(new_n396), .B2(KEYINPUT79), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT5), .ZN(new_n398));
  XOR2_X1   g197(.A(G1gat), .B(G29gat), .Z(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  AOI211_X1 g203(.A(new_n404), .B(new_n394), .C1(new_n395), .C2(new_n384), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n405), .A2(new_n406), .B1(new_n393), .B2(new_n391), .ZN(new_n407));
  AND4_X1   g206(.A1(KEYINPUT6), .A2(new_n398), .A3(new_n403), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n398), .A2(new_n407), .ZN(new_n409));
  INV_X1    g208(.A(new_n403), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n403), .A3(new_n407), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G226gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n203), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(KEYINPUT29), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n358), .A2(KEYINPUT74), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT74), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n332), .A2(new_n419), .A3(new_n346), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n358), .A2(new_n414), .A3(new_n203), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n236), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(new_n415), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n358), .A2(new_n416), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n235), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n423), .A2(new_n426), .ZN(new_n433));
  INV_X1    g232(.A(new_n429), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n426), .A4(new_n429), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n413), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n296), .A2(new_n382), .A3(new_n383), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n296), .A2(new_n383), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT70), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n379), .A2(new_n446), .A3(new_n381), .ZN(new_n447));
  INV_X1    g246(.A(new_n376), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n446), .B1(new_n379), .B2(new_n381), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n412), .B(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n408), .B1(new_n453), .B2(new_n411), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n454), .A2(KEYINPUT35), .A3(new_n437), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n445), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n442), .A2(new_n443), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n382), .A2(KEYINPUT36), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n451), .B2(KEYINPUT36), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n235), .B1(new_n421), .B2(new_n422), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n424), .A2(new_n236), .A3(new_n425), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT37), .A3(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT85), .Z(new_n463));
  OAI21_X1  g262(.A(new_n434), .B1(new_n433), .B2(KEYINPUT37), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT38), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n433), .A2(KEYINPUT37), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT38), .B1(new_n467), .B2(new_n464), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n466), .A2(new_n454), .A3(new_n430), .A4(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n391), .A2(new_n393), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n395), .A2(new_n394), .A3(new_n384), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n472), .B(new_n410), .C1(new_n470), .C2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT40), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n437), .A3(new_n453), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n445), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n444), .B1(new_n413), .B2(new_n437), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n482));
  INV_X1    g281(.A(G57gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G64gat), .ZN(new_n484));
  INV_X1    g283(.A(G64gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G57gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n488), .B2(new_n487), .ZN(new_n490));
  XOR2_X1   g289(.A(G71gat), .B(G78gat), .Z(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n482), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT94), .B1(new_n483), .B2(G64gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n486), .B1(new_n484), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT21), .ZN(new_n500));
  XNOR2_X1  g299(.A(G127gat), .B(G155gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n499), .A2(KEYINPUT21), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G8gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  AOI21_X1  g307(.A(G1gat), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n507), .B(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n502), .B(new_n511), .Z(new_n512));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT95), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G183gat), .B(G211gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n512), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G134gat), .B(G162gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  INV_X1    g326(.A(G85gat), .ZN(new_n528));
  INV_X1    g327(.A(G92gat), .ZN(new_n529));
  AOI22_X1  g328(.A1(KEYINPUT8), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n531), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT88), .Z(new_n536));
  NOR2_X1   g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n535), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT87), .A3(new_n542), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT87), .B1(new_n546), .B2(new_n542), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n534), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(KEYINPUT89), .A3(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT89), .B1(new_n550), .B2(new_n551), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n531), .A2(new_n533), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n531), .A2(new_n533), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n561), .A2(new_n550), .B1(KEYINPUT41), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n542), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n569), .A2(new_n547), .B1(new_n540), .B2(new_n544), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n570), .B2(KEYINPUT17), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n552), .B1(new_n571), .B2(new_n554), .ZN(new_n572));
  INV_X1    g371(.A(new_n564), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT98), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n522), .B1(new_n565), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT96), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n574), .A3(new_n522), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n575), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n561), .A2(new_n499), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n534), .A2(new_n498), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n561), .A2(new_n499), .A3(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G230gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n203), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G176gat), .B(G204gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  AND2_X1   g398(.A1(new_n587), .A2(new_n589), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n596), .B(new_n599), .C1(new_n600), .C2(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(new_n599), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n595), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n594), .B1(new_n590), .B2(new_n591), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n520), .A2(new_n586), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n510), .B1(KEYINPUT17), .B2(new_n570), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n555), .B2(new_n556), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n510), .A2(new_n550), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT18), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n611), .B(KEYINPUT13), .Z(new_n616));
  NOR2_X1   g415(.A1(new_n510), .A2(new_n550), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(KEYINPUT91), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n510), .A2(new_n621), .A3(new_n550), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n616), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n611), .A4(new_n612), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n615), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G197gat), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT11), .B(G169gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n615), .A2(new_n624), .A3(new_n633), .A4(new_n625), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n608), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n481), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n413), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g439(.A1(new_n481), .A2(new_n637), .ZN(new_n641));
  INV_X1    g440(.A(new_n437), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n648), .A2(G8gat), .B1(new_n643), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n649), .B1(new_n646), .B2(new_n647), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n437), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT99), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n650), .B1(new_n658), .B2(new_n645), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n653), .B1(new_n656), .B2(new_n660), .ZN(G1325gat));
  AOI21_X1  g460(.A(G15gat), .B1(new_n638), .B2(new_n451), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  INV_X1    g462(.A(new_n459), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n638), .A2(G15gat), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n641), .A2(new_n445), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  AOI21_X1  g468(.A(new_n586), .B1(new_n457), .B2(new_n480), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n413), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n520), .A2(new_n636), .A3(new_n606), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n671), .A2(G29gat), .A3(new_n672), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  AND2_X1   g475(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n582), .A2(new_n585), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n481), .B2(new_n680), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n586), .B(new_n677), .C1(new_n457), .C2(new_n480), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n673), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n672), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n676), .A2(new_n684), .ZN(G1328gat));
  NOR4_X1   g484(.A1(new_n671), .A2(G36gat), .A3(new_n642), .A4(new_n674), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT46), .ZN(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n683), .B2(new_n642), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1329gat));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n690));
  INV_X1    g489(.A(G43gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n451), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n683), .A2(new_n459), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1330gat));
  OAI211_X1 g495(.A(new_n444), .B(new_n673), .C1(new_n681), .C2(new_n682), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n445), .A2(G50gat), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n690), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT103), .B(KEYINPUT48), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n697), .A2(G50gat), .B1(new_n690), .B2(new_n699), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n701), .A2(new_n705), .ZN(G1331gat));
  NOR4_X1   g505(.A1(new_n680), .A2(new_n519), .A3(new_n635), .A4(new_n607), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n481), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n672), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT104), .B(G57gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  INV_X1    g510(.A(new_n708), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n437), .B(KEYINPUT105), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT106), .Z(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1333gat));
  OAI21_X1  g518(.A(G71gat), .B1(new_n708), .B2(new_n459), .ZN(new_n720));
  INV_X1    g519(.A(G71gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n451), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n708), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g523(.A1(new_n712), .A2(new_n444), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n520), .A2(new_n635), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n481), .A2(KEYINPUT51), .A3(new_n680), .A4(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n670), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n670), .A2(new_n727), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n732), .A2(KEYINPUT109), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n730), .A2(new_n736), .A3(new_n731), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n738), .A2(new_n528), .A3(new_n413), .A4(new_n606), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n520), .A2(new_n635), .A3(new_n607), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n681), .B2(new_n682), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g542(.A(KEYINPUT107), .B(new_n740), .C1(new_n681), .C2(new_n682), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n413), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G85gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n739), .A2(new_n746), .ZN(G1336gat));
  NAND3_X1  g546(.A1(new_n713), .A2(new_n529), .A3(new_n606), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n734), .A2(new_n733), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n732), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n743), .A2(new_n437), .A3(new_n744), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G92gat), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n748), .B1(new_n735), .B2(new_n737), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n741), .B2(new_n714), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n753), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n756), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n743), .A2(new_n664), .A3(new_n744), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n760), .A3(new_n664), .A4(new_n744), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(G99gat), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n607), .A2(G99gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n738), .A2(new_n451), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1338gat));
  OR3_X1    g564(.A1(new_n445), .A2(G106gat), .A3(new_n607), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n732), .B2(new_n749), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n444), .A3(new_n744), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(G106gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n735), .B2(new_n737), .ZN(new_n771));
  OAI21_X1  g570(.A(G106gat), .B1(new_n741), .B2(new_n445), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n770), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n773), .ZN(G1339gat));
  NOR3_X1   g573(.A1(new_n619), .A2(new_n616), .A3(new_n623), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n611), .B1(new_n610), .B2(new_n612), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n630), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n634), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n596), .A2(KEYINPUT54), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n599), .B1(new_n604), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n601), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT55), .B1(new_n780), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n680), .A2(new_n778), .A3(new_n786), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n635), .A2(new_n786), .B1(new_n778), .B2(new_n606), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n680), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n520), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n787), .B(KEYINPUT112), .C1(new_n788), .C2(new_n680), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT111), .B1(new_n608), .B2(new_n635), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n680), .A2(new_n519), .A3(new_n606), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n636), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n672), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n445), .A2(new_n382), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n714), .ZN(new_n801));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n635), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n635), .A2(new_n786), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n778), .A2(new_n606), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n680), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND4_X1   g604(.A1(new_n582), .A2(new_n786), .A3(new_n778), .A4(new_n585), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n790), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n519), .A3(new_n792), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n796), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n713), .A2(new_n672), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n451), .A2(new_n810), .A3(new_n445), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n636), .A2(new_n301), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(G1340gat));
  AOI21_X1  g613(.A(G120gat), .B1(new_n801), .B2(new_n606), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n607), .A2(new_n299), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n812), .B2(new_n816), .ZN(G1341gat));
  INV_X1    g616(.A(G127gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n818), .A3(new_n520), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n812), .A2(new_n520), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n818), .B2(new_n820), .ZN(G1342gat));
  AOI21_X1  g620(.A(G134gat), .B1(KEYINPUT113), .B2(KEYINPUT56), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n800), .A2(new_n642), .A3(new_n680), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n812), .A2(new_n680), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G134gat), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1343gat));
  AOI21_X1  g628(.A(new_n445), .B1(new_n808), .B2(new_n809), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n459), .A2(new_n811), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n789), .A2(new_n519), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n445), .B1(new_n809), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n832), .B(new_n833), .C1(new_n831), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G141gat), .B1(new_n836), .B2(new_n636), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n810), .A2(new_n413), .A3(new_n459), .A4(new_n444), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n713), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n635), .A2(new_n259), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT115), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT58), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n249), .A2(KEYINPUT59), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n836), .B2(new_n607), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n834), .B1(new_n635), .B2(new_n608), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n831), .A3(new_n444), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(new_n606), .C1(new_n830), .C2(new_n831), .ZN(new_n849));
  INV_X1    g648(.A(new_n833), .ZN(new_n850));
  OAI21_X1  g649(.A(G148gat), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT116), .B1(new_n851), .B2(KEYINPUT59), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n249), .A3(new_n606), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1345gat));
  OAI21_X1  g655(.A(G155gat), .B1(new_n836), .B2(new_n519), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n240), .A3(new_n520), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT117), .ZN(G1346gat));
  OAI21_X1  g659(.A(G162gat), .B1(new_n836), .B2(new_n586), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n680), .A2(new_n241), .A3(new_n642), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n838), .B2(new_n862), .ZN(G1347gat));
  NOR2_X1   g662(.A1(new_n797), .A2(new_n413), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n799), .A2(new_n713), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(G169gat), .B1(new_n866), .B2(new_n635), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n642), .A2(new_n413), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n451), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n810), .A2(new_n445), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n810), .A2(KEYINPUT118), .A3(new_n445), .A4(new_n869), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n636), .A2(new_n334), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n874), .B2(new_n875), .ZN(G1348gat));
  NAND3_X1  g675(.A1(new_n866), .A2(new_n335), .A3(new_n606), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n874), .A2(new_n606), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n335), .ZN(G1349gat));
  NAND3_X1  g678(.A1(new_n872), .A2(new_n520), .A3(new_n873), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G183gat), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n520), .A2(new_n339), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n864), .A2(KEYINPUT119), .A3(new_n865), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n810), .A2(new_n672), .A3(new_n865), .A4(new_n882), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(KEYINPUT121), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT60), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n880), .A2(G183gat), .B1(new_n883), .B2(new_n886), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT120), .B1(new_n891), .B2(KEYINPUT121), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT60), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n891), .B2(KEYINPUT120), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n892), .B2(new_n894), .ZN(G1350gat));
  AOI21_X1  g694(.A(new_n340), .B1(new_n874), .B2(new_n680), .ZN(new_n896));
  OR2_X1    g695(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g696(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n864), .A2(new_n340), .A3(new_n680), .A4(new_n865), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT122), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n899), .B(new_n901), .C1(new_n896), .C2(new_n897), .ZN(G1351gat));
  XOR2_X1   g701(.A(KEYINPUT124), .B(G197gat), .Z(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n797), .B2(new_n445), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n459), .A2(new_n868), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n848), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n907), .B2(new_n636), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n664), .A2(new_n445), .A3(new_n714), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n864), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n636), .A2(new_n903), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1352gat));
  OR3_X1    g711(.A1(new_n910), .A2(G204gat), .A3(new_n607), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G204gat), .B1(new_n849), .B2(new_n905), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n917), .B(new_n918), .C1(new_n915), .C2(new_n913), .ZN(G1353gat));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n520), .A3(new_n848), .A4(new_n906), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n520), .A2(new_n212), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n910), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n910), .B2(new_n924), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n920), .A2(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n922), .A2(new_n920), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n907), .B2(new_n586), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n680), .A2(new_n213), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n910), .B2(new_n932), .ZN(G1355gat));
endmodule


