//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT73), .A2(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT73), .A2(G125), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G140), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT74), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G140), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(KEYINPUT74), .A3(G140), .A4(new_n190), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n188), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT16), .A2(G140), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT73), .A2(G125), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT73), .A2(G125), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT75), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n204), .B(new_n199), .C1(new_n200), .C2(new_n201), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n187), .B1(new_n198), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n200), .A2(new_n201), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n194), .B1(new_n208), .B2(G140), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NOR4_X1   g024(.A1(new_n200), .A2(new_n201), .A3(new_n192), .A4(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT16), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n189), .A2(new_n190), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n204), .B1(new_n213), .B2(new_n199), .ZN(new_n214));
  INV_X1    g028(.A(new_n205), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(G146), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n207), .A2(new_n217), .A3(KEYINPUT76), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n219), .B(new_n187), .C1(new_n198), .C2(new_n206), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G128), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G110), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n222), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT24), .B(G110), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n218), .A2(new_n220), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G125), .B(G140), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n187), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n228), .A2(new_n229), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n231), .A2(new_n232), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n217), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT22), .B(G137), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n242), .B(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT72), .B(G902), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n235), .A2(new_n240), .A3(new_n245), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G217), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n248), .B2(G234), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(new_n249), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(G902), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n262), .B(KEYINPUT27), .Z(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT64), .B1(new_n267), .B2(G146), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n187), .A3(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n267), .A2(G146), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n274));
  OAI21_X1  g088(.A(G128), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G143), .B(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G137), .ZN(new_n283));
  INV_X1    g097(.A(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT11), .A3(G134), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(G137), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n283), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n282), .A2(G137), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n284), .A2(G134), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT65), .B(G131), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT65), .ZN(new_n292));
  XNOR2_X1  g106(.A(G134), .B(G137), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n280), .A2(new_n288), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G113), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G119), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n297), .B2(new_n298), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n283), .A2(new_n285), .A3(new_n287), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n288), .ZN(new_n308));
  AND2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NOR2_X1   g123(.A1(KEYINPUT0), .A2(G128), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n272), .A2(new_n311), .B1(new_n277), .B2(new_n309), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n295), .A2(new_n305), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n308), .A2(new_n312), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n294), .A2(new_n288), .A3(new_n291), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n272), .A2(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n317), .B(new_n320), .C1(new_n321), .C2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n295), .A2(new_n318), .A3(new_n319), .A4(new_n313), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n316), .B1(new_n327), .B2(new_n304), .ZN(new_n328));
  AOI211_X1 g142(.A(new_n315), .B(new_n305), .C1(new_n325), .C2(new_n326), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n266), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n304), .B1(new_n321), .B2(new_n324), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n314), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n314), .A2(new_n333), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n331), .A2(new_n332), .B1(new_n265), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n330), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT68), .B(new_n266), .C1(new_n328), .C2(new_n329), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(KEYINPUT31), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n348), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(new_n350), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n342), .B2(new_n346), .ZN(new_n355));
  INV_X1    g169(.A(G472), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n328), .A2(new_n329), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n265), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n337), .A2(new_n266), .A3(new_n339), .A4(new_n340), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n248), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n340), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n314), .A2(KEYINPUT71), .A3(new_n333), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n335), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n265), .A2(new_n359), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n362), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n356), .B1(new_n361), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n355), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n260), .B1(new_n351), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  INV_X1    g193(.A(G902), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n243), .A2(G227), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g198(.A(new_n308), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n187), .A2(G143), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n221), .B1(new_n386), .B2(KEYINPUT1), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n279), .B1(new_n387), .B2(new_n277), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G104), .ZN(new_n390));
  AND2_X1   g204(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(G104), .A3(new_n389), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G107), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n394), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n389), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(KEYINPUT80), .A3(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n399), .A2(new_n409), .A3(new_n402), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n399), .B2(new_n402), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n323), .A2(new_n404), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n407), .A2(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  INV_X1    g229(.A(new_n393), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n396), .A2(new_n398), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n415), .B(G101), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n312), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n401), .B1(new_n400), .B2(new_n395), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n394), .B1(new_n421), .B2(new_n393), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT79), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G101), .B1(new_n416), .B2(new_n417), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT4), .A4(new_n399), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n419), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n385), .B1(new_n414), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n411), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n399), .A2(new_n409), .A3(new_n402), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n413), .A3(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n403), .A2(KEYINPUT80), .A3(new_n404), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT80), .B1(new_n403), .B2(new_n404), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n435), .A2(new_n308), .A3(new_n427), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n384), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n399), .A2(new_n402), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n323), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n385), .B1(new_n439), .B2(new_n403), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n440), .A2(KEYINPUT12), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n403), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT12), .A3(new_n308), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n440), .A2(KEYINPUT12), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT82), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n407), .A2(new_n408), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n428), .A2(new_n449), .A3(new_n385), .A4(new_n432), .ZN(new_n450));
  INV_X1    g264(.A(new_n384), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n445), .A2(new_n448), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n362), .B1(new_n437), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n381), .B1(new_n453), .B2(new_n379), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n429), .B2(new_n436), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n441), .A2(new_n444), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT77), .B1(new_n450), .B2(new_n457), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n455), .A2(new_n458), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G469), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n378), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n423), .A2(new_n426), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n418), .A2(new_n304), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n225), .A2(G116), .ZN(new_n470));
  INV_X1    g284(.A(G116), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G119), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT5), .ZN(new_n473));
  OAI21_X1  g287(.A(G113), .B1(new_n470), .B2(KEYINPUT5), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n303), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n410), .A2(new_n411), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n466), .B1(new_n423), .B2(new_n426), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT83), .B1(new_n479), .B2(new_n476), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT84), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NOR4_X1   g297(.A1(new_n479), .A2(new_n476), .A3(KEYINPUT85), .A4(new_n482), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n485));
  INV_X1    g299(.A(new_n475), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n465), .A2(new_n467), .B1(new_n412), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n482), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n483), .B(KEYINPUT6), .C1(new_n484), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n312), .A2(new_n213), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n213), .B2(new_n323), .ZN(new_n492));
  INV_X1    g306(.A(G224), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(G953), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT87), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n492), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n497));
  NAND4_X1  g311(.A1(new_n478), .A2(new_n480), .A3(new_n482), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT7), .B1(new_n493), .B2(G953), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n492), .B(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n482), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n438), .A2(new_n475), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n399), .A2(KEYINPUT88), .A3(new_n402), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n475), .B1(new_n438), .B2(new_n504), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT89), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n438), .A2(new_n504), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n486), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n506), .A3(new_n505), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT89), .B1(new_n513), .B2(new_n503), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n501), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT90), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n468), .A2(new_n477), .A3(new_n488), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT85), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n487), .A2(new_n485), .A3(new_n488), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(new_n501), .C1(new_n510), .C2(new_n514), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G210), .B1(G237), .B2(G902), .ZN(new_n524));
  AND4_X1   g338(.A1(new_n380), .A2(new_n499), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n500), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n492), .B(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n530), .B2(new_n509), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n531), .A2(new_n521), .B1(new_n518), .B2(new_n519), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n532), .B2(new_n516), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n524), .B1(new_n533), .B2(new_n499), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n464), .B1(new_n525), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n463), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G475), .ZN(new_n537));
  INV_X1    g351(.A(G237), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n243), .A3(G214), .ZN(new_n539));
  AND2_X1   g353(.A1(KEYINPUT91), .A2(G143), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT91), .A2(G143), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n261), .B(G214), .C1(KEYINPUT91), .C2(G143), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT18), .A2(G131), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n196), .A2(G146), .A3(new_n197), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n237), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(KEYINPUT17), .A3(G131), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n544), .B(G131), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n218), .A2(new_n220), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n218), .A2(KEYINPUT95), .A3(new_n220), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G113), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT93), .B(G104), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(KEYINPUT97), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n558), .B2(new_n563), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n537), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n562), .B(new_n550), .C1(new_n556), .C2(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n217), .A2(new_n552), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n196), .A2(KEYINPUT19), .A3(new_n197), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT19), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n236), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n196), .A2(new_n571), .A3(KEYINPUT19), .A4(new_n197), .ZN(new_n575));
  AOI21_X1  g389(.A(G146), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n549), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n562), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n577), .B2(new_n562), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT96), .B1(new_n568), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n554), .A2(new_n555), .ZN(new_n585));
  INV_X1    g399(.A(new_n553), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n557), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n561), .A3(new_n549), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n577), .A2(new_n562), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n579), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(G475), .A2(G902), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n583), .A2(new_n584), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  AND4_X1   g409(.A1(new_n595), .A2(new_n592), .A3(new_n584), .A4(new_n593), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n567), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G952), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(G953), .ZN(new_n599));
  INV_X1    g413(.A(G234), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n538), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n243), .B(new_n248), .C1(G234), .C2(G237), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT21), .B(G898), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G478), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT15), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n267), .A2(G128), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n221), .A2(G143), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n282), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n471), .A2(KEYINPUT14), .A3(G122), .ZN(new_n613));
  XNOR2_X1  g427(.A(G116), .B(G122), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(G107), .B(new_n613), .C1(new_n615), .C2(KEYINPUT14), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n389), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n612), .A2(new_n620), .A3(new_n616), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n615), .A2(G107), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(new_n617), .B1(new_n282), .B2(new_n611), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n609), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n610), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n609), .A2(new_n624), .ZN(new_n627));
  OAI21_X1  g441(.A(G134), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n619), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n376), .A2(new_n253), .A3(G953), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT99), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n632), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(new_n619), .A3(new_n621), .A4(new_n629), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n362), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n608), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n248), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n638), .B1(new_n643), .B2(new_n608), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n597), .A2(new_n605), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n375), .A2(new_n536), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT101), .B(G101), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G3));
  AOI21_X1  g463(.A(new_n356), .B1(new_n347), .B2(new_n248), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n352), .B1(new_n342), .B2(new_n346), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n463), .A2(new_n650), .A3(new_n260), .A4(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n633), .B(new_n657), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n656), .A2(new_n658), .B1(new_n655), .B2(new_n639), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n362), .A2(new_n606), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n659), .A2(new_n660), .B1(new_n606), .B2(new_n640), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n597), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n605), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n464), .B(new_n664), .C1(new_n525), .C2(new_n534), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n652), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G104), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND3_X1  g484(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n558), .A2(new_n561), .B1(new_n590), .B2(new_n579), .ZN(new_n672));
  INV_X1    g486(.A(new_n593), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n584), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n645), .A2(new_n567), .A3(new_n671), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  XNOR2_X1  g493(.A(new_n241), .B(KEYINPUT105), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n246), .A2(KEYINPUT36), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(new_n258), .B1(new_n252), .B2(new_n254), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n650), .A2(new_n684), .A3(new_n651), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n536), .A3(new_n646), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AOI21_X1  g502(.A(new_n684), .B1(new_n351), .B2(new_n374), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n602), .B1(new_n603), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n675), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(new_n536), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  NAND2_X1  g508(.A1(new_n347), .A2(new_n353), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n266), .B1(new_n314), .B2(new_n334), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n344), .A2(new_n345), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n380), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G472), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n651), .A2(KEYINPUT32), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n464), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n683), .A2(new_n258), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n255), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n595), .B1(new_n588), .B2(new_n591), .ZN(new_n709));
  OAI22_X1  g523(.A1(new_n709), .A2(KEYINPUT20), .B1(new_n672), .B2(new_n673), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n592), .A2(new_n595), .A3(new_n584), .A4(new_n593), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n566), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n691), .B(KEYINPUT39), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n462), .A2(new_n713), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n712), .B(new_n644), .C1(new_n714), .C2(KEYINPUT40), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n716));
  INV_X1    g530(.A(new_n524), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n522), .A2(new_n520), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n531), .A2(new_n521), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n380), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n717), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n533), .A2(new_n499), .A3(new_n524), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n708), .A2(new_n715), .A3(new_n716), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  NOR3_X1   g543(.A1(new_n712), .A2(new_n661), .A3(new_n691), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n689), .A2(new_n536), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  NAND2_X1  g546(.A1(new_n437), .A2(new_n452), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n248), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n453), .A2(new_n379), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n377), .A3(new_n736), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n737), .B(new_n260), .C1(new_n351), .C2(new_n374), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n666), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  INV_X1    g554(.A(new_n260), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n735), .A2(new_n377), .A3(new_n736), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n355), .A2(new_n373), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n703), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n710), .A2(new_n711), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n661), .B1(new_n745), .B2(new_n567), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n705), .B1(new_n722), .B2(new_n723), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n664), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n739), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT41), .B(G113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G15));
  NAND2_X1  g566(.A1(new_n738), .A2(new_n676), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n535), .B2(new_n737), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n747), .A2(KEYINPUT109), .A3(new_n742), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n646), .A3(new_n689), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND4_X1  g574(.A1(new_n735), .A2(new_n377), .A3(new_n736), .A4(new_n664), .ZN(new_n761));
  INV_X1    g575(.A(new_n370), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n762), .A2(new_n265), .B1(new_n331), .B2(new_n332), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n352), .B1(new_n763), .B2(new_n346), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n260), .A2(new_n650), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n535), .A2(new_n712), .A3(new_n644), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  INV_X1    g582(.A(new_n691), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n746), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n712), .A2(new_n661), .A3(new_n771), .A4(new_n691), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n650), .A2(new_n684), .A3(new_n764), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n758), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  NAND3_X1  g590(.A1(new_n722), .A2(new_n464), .A3(new_n723), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n463), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n375), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n779), .A3(KEYINPUT42), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n597), .A2(new_n662), .A3(new_n769), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n771), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n746), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n375), .A2(new_n778), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  NAND3_X1  g603(.A1(new_n375), .A2(new_n778), .A3(new_n692), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  INV_X1    g605(.A(new_n777), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n707), .B1(new_n650), .B2(new_n651), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n712), .A2(new_n662), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT43), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT43), .B1(new_n712), .B2(new_n662), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n793), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n792), .B1(new_n799), .B2(KEYINPUT44), .ZN(new_n800));
  INV_X1    g614(.A(new_n793), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n801), .B(KEYINPUT44), .C1(new_n803), .C2(new_n797), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n460), .A2(KEYINPUT45), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n807));
  OAI221_X1 g621(.A(new_n807), .B1(new_n459), .B2(new_n451), .C1(new_n455), .C2(new_n458), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n806), .A2(G469), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n381), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT46), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n809), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n810), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n736), .A4(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n804), .A2(new_n816), .A3(new_n377), .A4(new_n713), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n800), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(KEYINPUT112), .B(G137), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G39));
  NOR2_X1   g634(.A1(new_n743), .A2(new_n703), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n260), .A3(new_n730), .A4(new_n792), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n377), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n816), .B2(new_n377), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND2_X1  g642(.A1(new_n735), .A2(new_n736), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT49), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n830), .A2(new_n705), .A3(new_n378), .A4(new_n260), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n724), .B(new_n725), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n704), .A3(new_n832), .A4(new_n795), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n378), .B(new_n691), .C1(new_n454), .C2(new_n461), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n836), .B(new_n684), .C1(new_n702), .C2(new_n703), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n747), .A2(new_n597), .A3(new_n645), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT114), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n347), .A2(new_n353), .B1(new_n700), .B2(G472), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n707), .B1(new_n351), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n766), .A2(new_n841), .A3(new_n842), .A4(new_n836), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n689), .B(new_n536), .C1(new_n692), .C2(new_n730), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n535), .A2(new_n755), .A3(new_n737), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT109), .B1(new_n747), .B2(new_n742), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n774), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(new_n848), .B2(new_n785), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n835), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n839), .A2(new_n843), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n775), .A3(KEYINPUT52), .A4(new_n845), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n738), .A2(new_n676), .B1(new_n765), .B2(new_n766), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n750), .A2(new_n759), .A3(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n566), .B(new_n644), .C1(new_n710), .C2(new_n711), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT113), .A3(new_n747), .A4(new_n664), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n712), .A2(new_n645), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n858), .B1(new_n859), .B2(new_n665), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n652), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n667), .A3(new_n647), .A4(new_n686), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n567), .A2(new_n644), .A3(new_n671), .A4(new_n674), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n689), .A2(new_n792), .A3(new_n836), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n774), .A2(new_n778), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n790), .B(new_n864), .C1(new_n785), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n855), .A2(new_n867), .A3(new_n788), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n834), .B1(new_n853), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n780), .A2(new_n787), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n750), .A2(new_n759), .A3(new_n854), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n852), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n862), .A2(new_n866), .A3(new_n834), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n759), .A2(new_n753), .A3(new_n767), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n788), .A3(KEYINPUT115), .A4(new_n750), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n869), .A2(new_n870), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT116), .ZN(new_n882));
  INV_X1    g696(.A(new_n868), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n883), .B2(new_n875), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n853), .A2(new_n868), .A3(new_n834), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n869), .A2(new_n887), .A3(new_n870), .A4(new_n880), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n777), .A2(new_n737), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n704), .A2(new_n889), .A3(new_n602), .A4(new_n741), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(new_n597), .A3(new_n662), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n601), .B1(new_n796), .B2(new_n798), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n889), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(new_n774), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n742), .A2(new_n705), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n727), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n650), .A2(new_n260), .A3(new_n764), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n892), .A2(new_n898), .A3(KEYINPUT50), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT50), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n602), .B(new_n899), .C1(new_n803), .C2(new_n797), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n832), .A2(new_n705), .A3(new_n742), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n896), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n829), .A2(new_n377), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n825), .A2(new_n826), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n902), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n792), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n895), .B(new_n905), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n758), .ZN(new_n911));
  OAI221_X1 g725(.A(new_n599), .B1(new_n890), .B2(new_n663), .C1(new_n902), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n375), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n893), .A2(KEYINPUT48), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT48), .B1(new_n893), .B2(new_n913), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n907), .A2(new_n909), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n900), .A2(new_n904), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(KEYINPUT117), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n895), .A4(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n917), .B1(new_n922), .B2(new_n896), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n882), .A2(new_n886), .A3(new_n888), .A4(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n598), .A2(new_n243), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n833), .B1(new_n926), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n243), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n869), .A2(new_n880), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n717), .A3(new_n362), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n490), .A2(new_n498), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n496), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT56), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n940), .B2(new_n933), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n942), .B2(new_n937), .ZN(G51));
  XNOR2_X1  g757(.A(new_n381), .B(KEYINPUT57), .ZN(new_n944));
  INV_X1    g758(.A(new_n881), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n870), .B1(new_n869), .B2(new_n880), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n733), .B(KEYINPUT120), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n932), .A2(new_n362), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(new_n809), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n930), .B1(new_n949), .B2(new_n951), .ZN(G54));
  NAND2_X1  g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n672), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n931), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n950), .A2(new_n672), .A3(new_n953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G60));
  NAND3_X1  g771(.A1(new_n882), .A2(new_n886), .A3(new_n888), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n659), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n659), .B(new_n961), .C1(new_n945), .C2(new_n946), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n931), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n964), .ZN(G63));
  AND2_X1   g779(.A1(new_n869), .A2(new_n880), .ZN(new_n966));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n256), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n869), .B2(new_n880), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n930), .B1(new_n970), .B2(new_n683), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT121), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT61), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n969), .B(new_n971), .C1(KEYINPUT121), .C2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n604), .B2(new_n493), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT122), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n873), .A2(new_n862), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(G953), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n935), .B1(G898), .B2(new_n243), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G69));
  NAND2_X1  g797(.A1(new_n690), .A2(G953), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n913), .A2(new_n838), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n816), .A3(new_n377), .A4(new_n713), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n827), .A2(new_n788), .A3(new_n790), .A4(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n800), .A2(new_n817), .ZN(new_n988));
  INV_X1    g802(.A(new_n849), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(KEYINPUT125), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT125), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n818), .B2(new_n849), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n987), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n984), .B1(new_n993), .B2(G953), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(KEYINPUT126), .B(new_n984), .C1(new_n993), .C2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n574), .A2(new_n575), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n327), .B(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n779), .B(new_n713), .C1(new_n746), .C2(new_n856), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n800), .B2(new_n817), .ZN(new_n1003));
  INV_X1    g817(.A(new_n826), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n822), .B1(new_n1004), .B2(new_n824), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n728), .A2(new_n775), .A3(new_n845), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n728), .A2(new_n775), .A3(new_n1009), .A4(new_n845), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT123), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1006), .B(new_n1008), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n1001), .B(new_n999), .C1(new_n1014), .C2(new_n243), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n988), .A2(new_n1008), .A3(new_n827), .A4(new_n1002), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n243), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n999), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT124), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n243), .B1(G227), .B2(G900), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1000), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1000), .B2(new_n1021), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n993), .B2(new_n980), .ZN(new_n1029));
  INV_X1    g843(.A(new_n357), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n265), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n931), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1032), .A2(KEYINPUT127), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1032), .A2(KEYINPUT127), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1014), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1028), .B1(new_n1035), .B2(new_n980), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1036), .A2(new_n265), .A3(new_n1030), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n884), .A2(new_n885), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n344), .A2(new_n345), .A3(new_n358), .ZN(new_n1039));
  NOR3_X1   g853(.A1(new_n1038), .A2(new_n1028), .A3(new_n1039), .ZN(new_n1040));
  NOR4_X1   g854(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .A4(new_n1040), .ZN(G57));
endmodule


