

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711;

  XNOR2_X1 U361 ( .A(n462), .B(n461), .ZN(n468) );
  OR2_X1 U362 ( .A1(n460), .A2(n479), .ZN(n462) );
  OR2_X1 U363 ( .A1(n632), .A2(n459), .ZN(n460) );
  INV_X2 U364 ( .A(n478), .ZN(n643) );
  XNOR2_X2 U365 ( .A(n355), .B(n354), .ZN(n520) );
  XNOR2_X1 U366 ( .A(n424), .B(KEYINPUT0), .ZN(n479) );
  XNOR2_X1 U367 ( .A(n450), .B(n345), .ZN(n404) );
  XNOR2_X1 U368 ( .A(n404), .B(n341), .ZN(n388) );
  INV_X1 U369 ( .A(G475), .ZN(n438) );
  XNOR2_X1 U370 ( .A(n353), .B(n352), .ZN(n666) );
  XNOR2_X1 U371 ( .A(n696), .B(n349), .ZN(n353) );
  XNOR2_X1 U372 ( .A(n511), .B(n510), .ZN(n512) );
  BUF_X1 U373 ( .A(n665), .Z(n674) );
  AND2_X1 U374 ( .A1(n574), .A2(G953), .ZN(n679) );
  XNOR2_X1 U375 ( .A(n388), .B(KEYINPUT93), .ZN(n696) );
  XNOR2_X1 U376 ( .A(n412), .B(n411), .ZN(n504) );
  NOR2_X1 U377 ( .A1(G902), .A2(n666), .ZN(n355) );
  XNOR2_X1 U378 ( .A(n552), .B(KEYINPUT83), .ZN(n553) );
  XNOR2_X1 U379 ( .A(n350), .B(G107), .ZN(n687) );
  XNOR2_X1 U380 ( .A(G104), .B(G110), .ZN(n350) );
  XNOR2_X1 U381 ( .A(n695), .B(n367), .ZN(n369) );
  XNOR2_X1 U382 ( .A(n366), .B(n365), .ZN(n367) );
  INV_X1 U383 ( .A(G143), .ZN(n343) );
  XNOR2_X1 U384 ( .A(n522), .B(KEYINPUT41), .ZN(n655) );
  NOR2_X1 U385 ( .A1(n632), .A2(n633), .ZN(n522) );
  XNOR2_X1 U386 ( .A(n455), .B(n454), .ZN(n495) );
  NOR2_X1 U387 ( .A1(n592), .A2(G902), .ZN(n390) );
  XNOR2_X1 U388 ( .A(n571), .B(n340), .ZN(n572) );
  BUF_X1 U389 ( .A(n495), .Z(n710) );
  XNOR2_X1 U390 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U391 ( .A(G122), .B(G131), .Z(n338) );
  XOR2_X1 U392 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n339) );
  XNOR2_X1 U393 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n340) );
  XOR2_X1 U394 ( .A(n347), .B(n346), .Z(n341) );
  XOR2_X1 U395 ( .A(n549), .B(KEYINPUT47), .Z(n342) );
  NAND2_X1 U396 ( .A1(n598), .A2(n486), .ZN(n492) );
  OR2_X1 U397 ( .A1(n492), .A2(n491), .ZN(n493) );
  NOR2_X1 U398 ( .A1(n618), .A2(n342), .ZN(n550) );
  XNOR2_X1 U399 ( .A(n348), .B(G140), .ZN(n349) );
  XNOR2_X1 U400 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U401 ( .A(n405), .B(n351), .ZN(n352) );
  NOR2_X1 U402 ( .A1(n471), .A2(n645), .ZN(n476) );
  XNOR2_X1 U403 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U404 ( .A(n439), .B(n438), .ZN(n482) );
  XNOR2_X1 U405 ( .A(n374), .B(n373), .ZN(n675) );
  XNOR2_X1 U406 ( .A(n666), .B(n667), .ZN(n668) );
  XNOR2_X1 U407 ( .A(n524), .B(KEYINPUT111), .ZN(n525) );
  BUF_X1 U408 ( .A(n504), .Z(n559) );
  XNOR2_X1 U409 ( .A(n526), .B(n525), .ZN(n709) );
  XNOR2_X2 U410 ( .A(G128), .B(KEYINPUT77), .ZN(n344) );
  XNOR2_X2 U411 ( .A(n344), .B(n343), .ZN(n450) );
  XNOR2_X1 U412 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n345) );
  XOR2_X1 U413 ( .A(KEYINPUT68), .B(G131), .Z(n347) );
  XNOR2_X1 U414 ( .A(G137), .B(G134), .ZN(n346) );
  INV_X1 U415 ( .A(G953), .ZN(n701) );
  AND2_X1 U416 ( .A1(G227), .A2(n701), .ZN(n348) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(G101), .ZN(n385) );
  XNOR2_X1 U418 ( .A(n687), .B(n385), .ZN(n405) );
  XNOR2_X1 U419 ( .A(G146), .B(KEYINPUT76), .ZN(n351) );
  XNOR2_X1 U420 ( .A(KEYINPUT70), .B(G469), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n520), .B(KEYINPUT1), .ZN(n471) );
  XNOR2_X1 U422 ( .A(KEYINPUT15), .B(G902), .ZN(n568) );
  NAND2_X1 U423 ( .A1(G234), .A2(n568), .ZN(n356) );
  XNOR2_X1 U424 ( .A(KEYINPUT20), .B(n356), .ZN(n375) );
  AND2_X1 U425 ( .A1(n375), .A2(G221), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n357), .B(KEYINPUT21), .ZN(n640) );
  INV_X1 U427 ( .A(G125), .ZN(n358) );
  NAND2_X1 U428 ( .A1(n358), .A2(G146), .ZN(n361) );
  INV_X1 U429 ( .A(G146), .ZN(n359) );
  NAND2_X1 U430 ( .A1(G125), .A2(n359), .ZN(n360) );
  NAND2_X1 U431 ( .A1(n361), .A2(n360), .ZN(n396) );
  XNOR2_X1 U432 ( .A(n396), .B(G140), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n362), .B(KEYINPUT10), .ZN(n695) );
  XOR2_X1 U434 ( .A(KEYINPUT81), .B(KEYINPUT94), .Z(n364) );
  XNOR2_X1 U435 ( .A(G137), .B(G110), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n364), .B(n363), .ZN(n366) );
  XOR2_X1 U437 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n365) );
  INV_X1 U438 ( .A(KEYINPUT24), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n374) );
  NAND2_X1 U440 ( .A1(G234), .A2(n701), .ZN(n370) );
  XOR2_X1 U441 ( .A(KEYINPUT8), .B(n370), .Z(n446) );
  NAND2_X1 U442 ( .A1(n446), .A2(G221), .ZN(n372) );
  XNOR2_X1 U443 ( .A(G119), .B(G128), .ZN(n371) );
  NOR2_X1 U444 ( .A1(n675), .A2(G902), .ZN(n379) );
  XOR2_X1 U445 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n377) );
  NAND2_X1 U446 ( .A1(G217), .A2(n375), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X2 U448 ( .A(n379), .B(n378), .ZN(n639) );
  NAND2_X1 U449 ( .A1(n640), .A2(n639), .ZN(n645) );
  XNOR2_X1 U450 ( .A(G472), .B(KEYINPUT71), .ZN(n391) );
  NOR2_X1 U451 ( .A1(G953), .A2(G237), .ZN(n430) );
  NAND2_X1 U452 ( .A1(n430), .A2(G210), .ZN(n381) );
  XOR2_X1 U453 ( .A(G146), .B(KEYINPUT73), .Z(n380) );
  XNOR2_X1 U454 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U455 ( .A(n382), .B(KEYINPUT5), .Z(n387) );
  XNOR2_X1 U456 ( .A(G116), .B(G113), .ZN(n384) );
  XNOR2_X1 U457 ( .A(KEYINPUT3), .B(G119), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n384), .B(n383), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n402), .B(n385), .ZN(n386) );
  XNOR2_X1 U460 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X1 U461 ( .A(n389), .B(n388), .ZN(n592) );
  XOR2_X1 U462 ( .A(n391), .B(n390), .Z(n478) );
  XNOR2_X1 U463 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n392) );
  XNOR2_X1 U464 ( .A(n478), .B(n392), .ZN(n538) );
  INV_X1 U465 ( .A(n538), .ZN(n393) );
  NAND2_X1 U466 ( .A1(n476), .A2(n393), .ZN(n395) );
  INV_X1 U467 ( .A(KEYINPUT33), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n395), .B(n394), .ZN(n625) );
  XOR2_X1 U469 ( .A(KEYINPUT18), .B(n396), .Z(n399) );
  NAND2_X1 U470 ( .A1(G224), .A2(n701), .ZN(n397) );
  XNOR2_X1 U471 ( .A(n397), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n399), .B(n398), .ZN(n403) );
  XNOR2_X1 U473 ( .A(KEYINPUT16), .B(G122), .ZN(n400) );
  XNOR2_X1 U474 ( .A(n400), .B(KEYINPUT72), .ZN(n401) );
  XNOR2_X1 U475 ( .A(n402), .B(n401), .ZN(n688) );
  XNOR2_X1 U476 ( .A(n403), .B(n688), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n407), .B(n406), .ZN(n582) );
  NAND2_X1 U479 ( .A1(n582), .A2(n568), .ZN(n412) );
  INV_X1 U480 ( .A(G902), .ZN(n409) );
  INV_X1 U481 ( .A(G237), .ZN(n408) );
  NAND2_X1 U482 ( .A1(n409), .A2(n408), .ZN(n413) );
  NAND2_X1 U483 ( .A1(n413), .A2(G210), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n410), .B(KEYINPUT78), .ZN(n411) );
  NAND2_X1 U485 ( .A1(n413), .A2(G214), .ZN(n629) );
  INV_X1 U486 ( .A(n629), .ZN(n414) );
  OR2_X1 U487 ( .A1(n504), .A2(n414), .ZN(n417) );
  XNOR2_X1 U488 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n415) );
  XNOR2_X1 U489 ( .A(n415), .B(KEYINPUT64), .ZN(n416) );
  XNOR2_X2 U490 ( .A(n417), .B(n416), .ZN(n546) );
  NAND2_X1 U491 ( .A1(G234), .A2(G237), .ZN(n418) );
  XNOR2_X1 U492 ( .A(n418), .B(KEYINPUT14), .ZN(n420) );
  NAND2_X1 U493 ( .A1(n420), .A2(G902), .ZN(n419) );
  XNOR2_X1 U494 ( .A(n419), .B(KEYINPUT92), .ZN(n505) );
  XNOR2_X1 U495 ( .A(G898), .B(KEYINPUT91), .ZN(n684) );
  NAND2_X1 U496 ( .A1(G953), .A2(n684), .ZN(n691) );
  OR2_X1 U497 ( .A1(n505), .A2(n691), .ZN(n422) );
  NAND2_X1 U498 ( .A1(G952), .A2(n420), .ZN(n661) );
  NOR2_X1 U499 ( .A1(n661), .A2(G953), .ZN(n509) );
  INV_X1 U500 ( .A(n509), .ZN(n421) );
  NAND2_X1 U501 ( .A1(n422), .A2(n421), .ZN(n423) );
  NAND2_X1 U502 ( .A1(n546), .A2(n423), .ZN(n424) );
  NOR2_X1 U503 ( .A1(n625), .A2(n479), .ZN(n425) );
  XNOR2_X1 U504 ( .A(n425), .B(KEYINPUT34), .ZN(n453) );
  XNOR2_X1 U505 ( .A(G113), .B(G143), .ZN(n426) );
  XNOR2_X1 U506 ( .A(n338), .B(n426), .ZN(n429) );
  XNOR2_X1 U507 ( .A(G104), .B(KEYINPUT96), .ZN(n427) );
  XNOR2_X1 U508 ( .A(n339), .B(n427), .ZN(n428) );
  XNOR2_X1 U509 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U510 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n432) );
  NAND2_X1 U511 ( .A1(G214), .A2(n430), .ZN(n431) );
  XNOR2_X1 U512 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U513 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U514 ( .A(n435), .B(n695), .ZN(n571) );
  NOR2_X1 U515 ( .A1(G902), .A2(n571), .ZN(n437) );
  XNOR2_X1 U516 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n436) );
  XNOR2_X1 U517 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U518 ( .A(G107), .B(G122), .Z(n441) );
  XNOR2_X1 U519 ( .A(G116), .B(G134), .ZN(n440) );
  XNOR2_X1 U520 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U521 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n443) );
  XNOR2_X1 U522 ( .A(KEYINPUT9), .B(KEYINPUT101), .ZN(n442) );
  XNOR2_X1 U523 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U524 ( .A(n445), .B(n444), .Z(n448) );
  NAND2_X1 U525 ( .A1(G217), .A2(n446), .ZN(n447) );
  XNOR2_X1 U526 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U527 ( .A(n450), .B(n449), .ZN(n671) );
  NOR2_X1 U528 ( .A1(G902), .A2(n671), .ZN(n451) );
  XOR2_X1 U529 ( .A(G478), .B(n451), .Z(n483) );
  NAND2_X1 U530 ( .A1(n482), .A2(n483), .ZN(n530) );
  INV_X1 U531 ( .A(n530), .ZN(n452) );
  NAND2_X1 U532 ( .A1(n453), .A2(n452), .ZN(n455) );
  INV_X1 U533 ( .A(KEYINPUT35), .ZN(n454) );
  NOR2_X1 U534 ( .A1(n495), .A2(KEYINPUT85), .ZN(n465) );
  NOR2_X1 U535 ( .A1(n639), .A2(n643), .ZN(n456) );
  AND2_X1 U536 ( .A1(n471), .A2(n456), .ZN(n463) );
  NOR2_X1 U537 ( .A1(n482), .A2(n483), .ZN(n458) );
  INV_X1 U538 ( .A(KEYINPUT104), .ZN(n457) );
  XNOR2_X1 U539 ( .A(n458), .B(n457), .ZN(n632) );
  INV_X1 U540 ( .A(n640), .ZN(n459) );
  INV_X1 U541 ( .A(KEYINPUT22), .ZN(n461) );
  AND2_X1 U542 ( .A1(n463), .A2(n468), .ZN(n605) );
  INV_X1 U543 ( .A(KEYINPUT44), .ZN(n490) );
  OR2_X1 U544 ( .A1(n605), .A2(n490), .ZN(n464) );
  NOR2_X1 U545 ( .A1(n465), .A2(n464), .ZN(n489) );
  BUF_X1 U546 ( .A(n471), .Z(n646) );
  NOR2_X1 U547 ( .A1(n646), .A2(n639), .ZN(n467) );
  INV_X1 U548 ( .A(KEYINPUT105), .ZN(n466) );
  XNOR2_X1 U549 ( .A(n467), .B(n466), .ZN(n469) );
  AND2_X2 U550 ( .A1(n468), .A2(n538), .ZN(n472) );
  NAND2_X1 U551 ( .A1(n469), .A2(n472), .ZN(n470) );
  XNOR2_X1 U552 ( .A(n470), .B(KEYINPUT32), .ZN(n588) );
  NAND2_X1 U553 ( .A1(n472), .A2(n471), .ZN(n474) );
  INV_X1 U554 ( .A(KEYINPUT84), .ZN(n473) );
  XNOR2_X1 U555 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U556 ( .A1(n475), .A2(n639), .ZN(n598) );
  NAND2_X1 U557 ( .A1(n643), .A2(n476), .ZN(n652) );
  NOR2_X1 U558 ( .A1(n652), .A2(n479), .ZN(n477) );
  XNOR2_X1 U559 ( .A(n477), .B(KEYINPUT31), .ZN(n615) );
  NOR2_X1 U560 ( .A1(n520), .A2(n645), .ZN(n529) );
  AND2_X1 U561 ( .A1(n529), .A2(n478), .ZN(n481) );
  INV_X1 U562 ( .A(n479), .ZN(n480) );
  NAND2_X1 U563 ( .A1(n481), .A2(n480), .ZN(n601) );
  NAND2_X1 U564 ( .A1(n615), .A2(n601), .ZN(n485) );
  XOR2_X1 U565 ( .A(KEYINPUT100), .B(n482), .Z(n484) );
  OR2_X1 U566 ( .A1(n484), .A2(n483), .ZN(n613) );
  NAND2_X1 U567 ( .A1(n484), .A2(n483), .ZN(n616) );
  NAND2_X1 U568 ( .A1(n613), .A2(n616), .ZN(n548) );
  NAND2_X1 U569 ( .A1(n485), .A2(n548), .ZN(n486) );
  INV_X1 U570 ( .A(n492), .ZN(n487) );
  AND2_X1 U571 ( .A1(n588), .A2(n487), .ZN(n488) );
  NAND2_X1 U572 ( .A1(n489), .A2(n488), .ZN(n494) );
  INV_X1 U573 ( .A(KEYINPUT85), .ZN(n497) );
  NAND2_X1 U574 ( .A1(n497), .A2(n490), .ZN(n491) );
  NAND2_X1 U575 ( .A1(n494), .A2(n493), .ZN(n501) );
  NOR2_X1 U576 ( .A1(n605), .A2(KEYINPUT44), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n588), .A2(n496), .ZN(n498) );
  NAND2_X1 U578 ( .A1(n498), .A2(n497), .ZN(n499) );
  NAND2_X1 U579 ( .A1(n710), .A2(n499), .ZN(n500) );
  NAND2_X1 U580 ( .A1(n501), .A2(n500), .ZN(n503) );
  XNOR2_X1 U581 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n502) );
  XNOR2_X2 U582 ( .A(n503), .B(n502), .ZN(n680) );
  XNOR2_X1 U583 ( .A(KEYINPUT38), .B(n559), .ZN(n630) );
  OR2_X1 U584 ( .A1(n701), .A2(n505), .ZN(n506) );
  NOR2_X1 U585 ( .A1(G900), .A2(n506), .ZN(n507) );
  XNOR2_X1 U586 ( .A(n507), .B(KEYINPUT106), .ZN(n508) );
  NOR2_X1 U587 ( .A1(n509), .A2(n508), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n629), .A2(n643), .ZN(n511) );
  NOR2_X1 U589 ( .A1(n536), .A2(n512), .ZN(n528) );
  AND2_X1 U590 ( .A1(n630), .A2(n528), .ZN(n513) );
  AND2_X1 U591 ( .A1(n513), .A2(n529), .ZN(n514) );
  XNOR2_X1 U592 ( .A(n514), .B(KEYINPUT39), .ZN(n555) );
  NOR2_X1 U593 ( .A1(n555), .A2(n613), .ZN(n516) );
  XNOR2_X1 U594 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n515) );
  XNOR2_X1 U595 ( .A(n516), .B(n515), .ZN(n711) );
  NAND2_X1 U596 ( .A1(n643), .A2(n640), .ZN(n517) );
  OR2_X1 U597 ( .A1(n536), .A2(n517), .ZN(n518) );
  NOR2_X1 U598 ( .A1(n639), .A2(n518), .ZN(n519) );
  XOR2_X1 U599 ( .A(KEYINPUT28), .B(n519), .Z(n521) );
  NOR2_X1 U600 ( .A1(n521), .A2(n520), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n630), .A2(n629), .ZN(n633) );
  INV_X1 U602 ( .A(n655), .ZN(n523) );
  NAND2_X1 U603 ( .A1(n547), .A2(n523), .ZN(n526) );
  XOR2_X1 U604 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n524) );
  NAND2_X1 U605 ( .A1(n711), .A2(n709), .ZN(n527) );
  XNOR2_X1 U606 ( .A(n527), .B(KEYINPUT46), .ZN(n534) );
  NAND2_X1 U607 ( .A1(n529), .A2(n528), .ZN(n531) );
  OR2_X1 U608 ( .A1(n531), .A2(n530), .ZN(n532) );
  OR2_X1 U609 ( .A1(n559), .A2(n532), .ZN(n587) );
  INV_X1 U610 ( .A(n587), .ZN(n533) );
  NOR2_X1 U611 ( .A1(n534), .A2(n533), .ZN(n551) );
  XOR2_X1 U612 ( .A(KEYINPUT86), .B(KEYINPUT112), .Z(n535) );
  XNOR2_X1 U613 ( .A(KEYINPUT36), .B(n535), .ZN(n544) );
  NOR2_X1 U614 ( .A1(n536), .A2(n639), .ZN(n537) );
  NAND2_X1 U615 ( .A1(n537), .A2(n640), .ZN(n539) );
  NOR2_X1 U616 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U617 ( .A1(n540), .A2(n629), .ZN(n541) );
  NOR2_X1 U618 ( .A1(n613), .A2(n541), .ZN(n556) );
  INV_X1 U619 ( .A(n559), .ZN(n542) );
  NAND2_X1 U620 ( .A1(n556), .A2(n542), .ZN(n543) );
  XOR2_X1 U621 ( .A(n544), .B(n543), .Z(n545) );
  NOR2_X1 U622 ( .A1(n646), .A2(n545), .ZN(n618) );
  NAND2_X1 U623 ( .A1(n547), .A2(n546), .ZN(n611) );
  INV_X1 U624 ( .A(n548), .ZN(n634) );
  NOR2_X1 U625 ( .A1(n611), .A2(n634), .ZN(n549) );
  AND2_X1 U626 ( .A1(n551), .A2(n550), .ZN(n554) );
  XNOR2_X1 U627 ( .A(KEYINPUT48), .B(KEYINPUT69), .ZN(n552) );
  XNOR2_X1 U628 ( .A(n554), .B(n553), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n555), .A2(n616), .ZN(n621) );
  XOR2_X1 U630 ( .A(KEYINPUT107), .B(n556), .Z(n557) );
  NAND2_X1 U631 ( .A1(n557), .A2(n646), .ZN(n558) );
  XNOR2_X1 U632 ( .A(KEYINPUT43), .B(n558), .ZN(n560) );
  AND2_X1 U633 ( .A1(n560), .A2(n559), .ZN(n590) );
  NOR2_X1 U634 ( .A1(n621), .A2(n590), .ZN(n561) );
  NAND2_X1 U635 ( .A1(n562), .A2(n561), .ZN(n698) );
  INV_X1 U636 ( .A(n698), .ZN(n563) );
  NAND2_X1 U637 ( .A1(n680), .A2(n563), .ZN(n565) );
  INV_X1 U638 ( .A(KEYINPUT2), .ZN(n564) );
  NAND2_X1 U639 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U640 ( .A(n566), .ZN(n622) );
  NOR2_X1 U641 ( .A1(n698), .A2(n564), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n680), .A2(n567), .ZN(n623) );
  INV_X1 U643 ( .A(n568), .ZN(n569) );
  NAND2_X1 U644 ( .A1(n623), .A2(n569), .ZN(n570) );
  NOR2_X4 U645 ( .A1(n622), .A2(n570), .ZN(n665) );
  NAND2_X1 U646 ( .A1(n665), .A2(G475), .ZN(n573) );
  XNOR2_X1 U647 ( .A(n573), .B(n572), .ZN(n575) );
  INV_X1 U648 ( .A(G952), .ZN(n574) );
  NOR2_X2 U649 ( .A1(n575), .A2(n679), .ZN(n577) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT65), .Z(n576) );
  XNOR2_X1 U651 ( .A(n577), .B(n576), .ZN(G60) );
  NAND2_X1 U652 ( .A1(n665), .A2(G210), .ZN(n584) );
  XNOR2_X1 U653 ( .A(KEYINPUT80), .B(KEYINPUT87), .ZN(n578) );
  XNOR2_X1 U654 ( .A(n578), .B(KEYINPUT55), .ZN(n579) );
  XNOR2_X1 U655 ( .A(KEYINPUT122), .B(n579), .ZN(n580) );
  XOR2_X1 U656 ( .A(n580), .B(KEYINPUT54), .Z(n581) );
  XNOR2_X1 U657 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X2 U659 ( .A1(n585), .A2(n679), .ZN(n586) );
  XNOR2_X1 U660 ( .A(n586), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U661 ( .A(n587), .B(G143), .ZN(G45) );
  XNOR2_X1 U662 ( .A(n588), .B(G119), .ZN(G21) );
  XNOR2_X1 U663 ( .A(G140), .B(KEYINPUT118), .ZN(n589) );
  XOR2_X1 U664 ( .A(n590), .B(n589), .Z(G42) );
  NAND2_X1 U665 ( .A1(n665), .A2(G472), .ZN(n594) );
  XNOR2_X1 U666 ( .A(KEYINPUT88), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U668 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X2 U669 ( .A1(n595), .A2(n679), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n596) );
  XNOR2_X1 U671 ( .A(n597), .B(n596), .ZN(G57) );
  XNOR2_X1 U672 ( .A(G101), .B(n598), .ZN(G3) );
  NOR2_X1 U673 ( .A1(n613), .A2(n601), .ZN(n600) );
  XNOR2_X1 U674 ( .A(G104), .B(KEYINPUT113), .ZN(n599) );
  XNOR2_X1 U675 ( .A(n600), .B(n599), .ZN(G6) );
  NOR2_X1 U676 ( .A1(n616), .A2(n601), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(G107), .B(n604), .ZN(G9) );
  XOR2_X1 U680 ( .A(G110), .B(n605), .Z(n606) );
  XNOR2_X1 U681 ( .A(KEYINPUT114), .B(n606), .ZN(G12) );
  NOR2_X1 U682 ( .A1(n611), .A2(n616), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n608) );
  XNOR2_X1 U684 ( .A(G128), .B(KEYINPUT116), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n610), .B(n609), .ZN(G30) );
  NOR2_X1 U687 ( .A1(n611), .A2(n613), .ZN(n612) );
  XOR2_X1 U688 ( .A(G146), .B(n612), .Z(G48) );
  NOR2_X1 U689 ( .A1(n613), .A2(n615), .ZN(n614) );
  XOR2_X1 U690 ( .A(G113), .B(n614), .Z(G15) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U692 ( .A(G116), .B(n617), .Z(G18) );
  XOR2_X1 U693 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n620) );
  XNOR2_X1 U694 ( .A(G125), .B(n618), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n620), .B(n619), .ZN(G27) );
  XOR2_X1 U696 ( .A(G134), .B(n621), .Z(G36) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT79), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n628) );
  BUF_X1 U699 ( .A(n625), .Z(n637) );
  NOR2_X1 U700 ( .A1(n655), .A2(n637), .ZN(n626) );
  NOR2_X1 U701 ( .A1(G953), .A2(n626), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n663) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n636) );
  NOR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n638) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n657) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U709 ( .A(KEYINPUT49), .B(n641), .Z(n642) );
  NOR2_X1 U710 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U711 ( .A(KEYINPUT119), .B(n644), .Z(n650) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n647), .B(KEYINPUT50), .ZN(n648) );
  XNOR2_X1 U714 ( .A(KEYINPUT120), .B(n648), .ZN(n649) );
  NAND2_X1 U715 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U716 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U717 ( .A(KEYINPUT51), .B(n653), .ZN(n654) );
  NOR2_X1 U718 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U719 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U720 ( .A(n658), .B(KEYINPUT52), .Z(n659) );
  XNOR2_X1 U721 ( .A(KEYINPUT121), .B(n659), .ZN(n660) );
  NOR2_X1 U722 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U723 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U724 ( .A(n664), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U725 ( .A1(n674), .A2(G469), .ZN(n669) );
  XOR2_X1 U726 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n667) );
  NOR2_X1 U727 ( .A1(n679), .A2(n670), .ZN(G54) );
  NAND2_X1 U728 ( .A1(n674), .A2(G478), .ZN(n672) );
  XNOR2_X1 U729 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U730 ( .A1(n679), .A2(n673), .ZN(G63) );
  NAND2_X1 U731 ( .A1(n674), .A2(G217), .ZN(n677) );
  XOR2_X1 U732 ( .A(n675), .B(KEYINPUT123), .Z(n676) );
  XNOR2_X1 U733 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U734 ( .A1(n679), .A2(n678), .ZN(G66) );
  INV_X1 U735 ( .A(n680), .ZN(n681) );
  NOR2_X1 U736 ( .A1(n681), .A2(G953), .ZN(n686) );
  NAND2_X1 U737 ( .A1(G953), .A2(G224), .ZN(n682) );
  XOR2_X1 U738 ( .A(KEYINPUT61), .B(n682), .Z(n683) );
  NOR2_X1 U739 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U740 ( .A1(n686), .A2(n685), .ZN(n693) );
  XNOR2_X1 U741 ( .A(n687), .B(G101), .ZN(n689) );
  XOR2_X1 U742 ( .A(n689), .B(n688), .Z(n690) );
  NAND2_X1 U743 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U744 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U745 ( .A(KEYINPUT124), .B(n694), .ZN(G69) );
  XOR2_X1 U746 ( .A(n696), .B(n695), .Z(n703) );
  INV_X1 U747 ( .A(n703), .ZN(n697) );
  XOR2_X1 U748 ( .A(n697), .B(KEYINPUT125), .Z(n699) );
  XNOR2_X1 U749 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U750 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U751 ( .A(KEYINPUT126), .B(n702), .ZN(n708) );
  XOR2_X1 U752 ( .A(G227), .B(n703), .Z(n704) );
  NAND2_X1 U753 ( .A1(n704), .A2(G900), .ZN(n705) );
  NAND2_X1 U754 ( .A1(G953), .A2(n705), .ZN(n706) );
  XOR2_X1 U755 ( .A(KEYINPUT127), .B(n706), .Z(n707) );
  NAND2_X1 U756 ( .A1(n708), .A2(n707), .ZN(G72) );
  XNOR2_X1 U757 ( .A(n709), .B(G137), .ZN(G39) );
  XNOR2_X1 U758 ( .A(G122), .B(n710), .ZN(G24) );
  XNOR2_X1 U759 ( .A(n711), .B(G131), .ZN(G33) );
endmodule

