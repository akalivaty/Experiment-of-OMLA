

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XNOR2_X1 U323 ( .A(KEYINPUT120), .B(n442), .ZN(n561) );
  XNOR2_X1 U324 ( .A(n343), .B(n342), .ZN(n550) );
  XNOR2_X1 U325 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U326 ( .A(n330), .B(n329), .ZN(n334) );
  NOR2_X1 U327 ( .A1(n508), .A2(n422), .ZN(n564) );
  XNOR2_X1 U328 ( .A(n341), .B(n340), .ZN(n342) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n443) );
  XOR2_X1 U330 ( .A(n440), .B(n439), .Z(n522) );
  XOR2_X1 U331 ( .A(n460), .B(KEYINPUT28), .Z(n524) );
  XNOR2_X1 U332 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U333 ( .A(n446), .B(n445), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G50GAT), .B(G162GAT), .Z(n326) );
  XOR2_X1 U335 ( .A(G78GAT), .B(G106GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G22GAT), .B(G218GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(n326), .B(n293), .Z(n295) );
  NAND2_X1 U339 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U341 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n297) );
  XNOR2_X1 U342 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n299), .B(n298), .Z(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT3), .B(G155GAT), .Z(n301) );
  XNOR2_X1 U346 ( .A(KEYINPUT2), .B(G148GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U348 ( .A(G141GAT), .B(n302), .Z(n324) );
  XNOR2_X1 U349 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n303), .B(KEYINPUT86), .ZN(n304) );
  XOR2_X1 U351 ( .A(n304), .B(KEYINPUT21), .Z(n306) );
  XNOR2_X1 U352 ( .A(G197GAT), .B(G204GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n409) );
  XNOR2_X1 U354 ( .A(n324), .B(n409), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n460) );
  XOR2_X1 U356 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n310) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(n311), .B(KEYINPUT5), .Z(n316) );
  XOR2_X1 U360 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n313) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n432) );
  XNOR2_X1 U363 ( .A(G29GAT), .B(G134GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n314), .B(G85GAT), .ZN(n337) );
  XNOR2_X1 U365 ( .A(n432), .B(n337), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U367 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n318) );
  XOR2_X1 U368 ( .A(G120GAT), .B(G57GAT), .Z(n391) );
  XOR2_X1 U369 ( .A(G1GAT), .B(G127GAT), .Z(n353) );
  XNOR2_X1 U370 ( .A(n391), .B(n353), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U372 ( .A(n320), .B(n319), .Z(n322) );
  XNOR2_X1 U373 ( .A(G162GAT), .B(KEYINPUT4), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n464) );
  XNOR2_X1 U376 ( .A(KEYINPUT91), .B(n464), .ZN(n508) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(G218GAT), .ZN(n416) );
  XNOR2_X1 U379 ( .A(n416), .B(n326), .ZN(n330) );
  AND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n328) );
  INV_X1 U381 ( .A(KEYINPUT64), .ZN(n327) );
  XOR2_X1 U382 ( .A(G43GAT), .B(KEYINPUT8), .Z(n332) );
  XNOR2_X1 U383 ( .A(KEYINPUT7), .B(KEYINPUT67), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n369) );
  XNOR2_X1 U385 ( .A(n369), .B(KEYINPUT11), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n343) );
  XOR2_X1 U387 ( .A(KEYINPUT70), .B(G92GAT), .Z(n336) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n384) );
  XNOR2_X1 U390 ( .A(n337), .B(n384), .ZN(n341) );
  XOR2_X1 U391 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n339) );
  XNOR2_X1 U392 ( .A(KEYINPUT73), .B(KEYINPUT9), .ZN(n338) );
  XOR2_X1 U393 ( .A(n339), .B(n338), .Z(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n345) );
  XNOR2_X1 U395 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U397 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n347) );
  XNOR2_X1 U398 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n361) );
  XOR2_X1 U401 ( .A(G64GAT), .B(G57GAT), .Z(n351) );
  XNOR2_X1 U402 ( .A(G155GAT), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n357) );
  XNOR2_X1 U404 ( .A(G71GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n352), .B(KEYINPUT13), .ZN(n383) );
  XOR2_X1 U406 ( .A(n383), .B(n353), .Z(n355) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U409 ( .A(n357), .B(n356), .Z(n359) );
  XOR2_X1 U410 ( .A(G15GAT), .B(G22GAT), .Z(n365) );
  XOR2_X1 U411 ( .A(G8GAT), .B(G183GAT), .Z(n405) );
  XNOR2_X1 U412 ( .A(n365), .B(n405), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n573) );
  XOR2_X1 U415 ( .A(G36GAT), .B(G50GAT), .Z(n363) );
  XNOR2_X1 U416 ( .A(G169GAT), .B(G29GAT), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U418 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U421 ( .A(n368), .B(KEYINPUT29), .Z(n371) );
  XNOR2_X1 U422 ( .A(n369), .B(KEYINPUT65), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n371), .B(n370), .ZN(n379) );
  XOR2_X1 U424 ( .A(G1GAT), .B(G197GAT), .Z(n373) );
  XNOR2_X1 U425 ( .A(G113GAT), .B(G141GAT), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U427 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n375) );
  XNOR2_X1 U428 ( .A(G8GAT), .B(KEYINPUT66), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U430 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n565) );
  XOR2_X1 U432 ( .A(KEYINPUT32), .B(KEYINPUT69), .Z(n381) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U435 ( .A(n382), .B(KEYINPUT33), .Z(n386) );
  XNOR2_X1 U436 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U438 ( .A(KEYINPUT31), .B(G85GAT), .Z(n388) );
  XNOR2_X1 U439 ( .A(G148GAT), .B(G204GAT), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U441 ( .A(n390), .B(n389), .Z(n393) );
  XOR2_X1 U442 ( .A(G176GAT), .B(G64GAT), .Z(n404) );
  XNOR2_X1 U443 ( .A(n391), .B(n404), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n570) );
  XNOR2_X1 U445 ( .A(n570), .B(KEYINPUT41), .ZN(n554) );
  NOR2_X1 U446 ( .A1(n565), .A2(n554), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n394), .B(KEYINPUT46), .ZN(n395) );
  NOR2_X1 U448 ( .A1(n573), .A2(n395), .ZN(n396) );
  NAND2_X1 U449 ( .A1(n550), .A2(n396), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n397), .B(KEYINPUT47), .ZN(n402) );
  XNOR2_X1 U451 ( .A(KEYINPUT74), .B(n550), .ZN(n535) );
  XNOR2_X1 U452 ( .A(KEYINPUT36), .B(n535), .ZN(n578) );
  INV_X1 U453 ( .A(n573), .ZN(n560) );
  NOR2_X1 U454 ( .A1(n578), .A2(n560), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n398), .B(KEYINPUT45), .ZN(n399) );
  NAND2_X1 U456 ( .A1(n399), .A2(n565), .ZN(n400) );
  NOR2_X1 U457 ( .A1(n400), .A2(n570), .ZN(n401) );
  NOR2_X1 U458 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n403), .B(KEYINPUT48), .ZN(n520) );
  XOR2_X1 U460 ( .A(KEYINPUT94), .B(G92GAT), .Z(n407) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U463 ( .A(n409), .B(n408), .Z(n411) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n420) );
  XOR2_X1 U466 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n418) );
  XNOR2_X1 U467 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n412), .B(KEYINPUT84), .ZN(n413) );
  XOR2_X1 U469 ( .A(n413), .B(KEYINPUT83), .Z(n415) );
  XNOR2_X1 U470 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n436) );
  XNOR2_X1 U472 ( .A(n436), .B(n416), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U474 ( .A(n420), .B(n419), .Z(n458) );
  NOR2_X1 U475 ( .A1(n520), .A2(n458), .ZN(n421) );
  XOR2_X1 U476 ( .A(KEYINPUT54), .B(n421), .Z(n422) );
  NAND2_X1 U477 ( .A1(n460), .A2(n564), .ZN(n423) );
  XNOR2_X1 U478 ( .A(KEYINPUT55), .B(n423), .ZN(n441) );
  XOR2_X1 U479 ( .A(G176GAT), .B(KEYINPUT82), .Z(n425) );
  XNOR2_X1 U480 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n440) );
  XOR2_X1 U482 ( .A(G190GAT), .B(G134GAT), .Z(n427) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G99GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U485 ( .A(G127GAT), .B(G183GAT), .Z(n429) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(G120GAT), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n438) );
  XOR2_X1 U489 ( .A(n432), .B(G71GAT), .Z(n434) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U494 ( .A1(n441), .A2(n522), .ZN(n442) );
  NOR2_X1 U495 ( .A1(n561), .A2(n535), .ZN(n446) );
  XNOR2_X1 U496 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n444) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n447), .B(KEYINPUT34), .ZN(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT98), .B(n448), .Z(n470) );
  NOR2_X1 U500 ( .A1(n565), .A2(n570), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n449), .B(KEYINPUT71), .ZN(n482) );
  NAND2_X1 U502 ( .A1(n573), .A2(n535), .ZN(n450) );
  XOR2_X1 U503 ( .A(KEYINPUT16), .B(n450), .Z(n468) );
  XOR2_X1 U504 ( .A(n458), .B(KEYINPUT27), .Z(n457) );
  NAND2_X1 U505 ( .A1(n457), .A2(n508), .ZN(n451) );
  XOR2_X1 U506 ( .A(KEYINPUT95), .B(n451), .Z(n519) );
  NOR2_X1 U507 ( .A1(n524), .A2(n519), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT96), .ZN(n454) );
  INV_X1 U509 ( .A(n522), .ZN(n453) );
  NAND2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n467) );
  NOR2_X1 U511 ( .A1(n522), .A2(n460), .ZN(n455) );
  XOR2_X1 U512 ( .A(KEYINPUT97), .B(n455), .Z(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT26), .B(n456), .ZN(n563) );
  NAND2_X1 U514 ( .A1(n563), .A2(n457), .ZN(n463) );
  INV_X1 U515 ( .A(n458), .ZN(n510) );
  NAND2_X1 U516 ( .A1(n522), .A2(n510), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n461), .Z(n462) );
  NAND2_X1 U519 ( .A1(n463), .A2(n462), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n477) );
  NAND2_X1 U522 ( .A1(n468), .A2(n477), .ZN(n495) );
  NOR2_X1 U523 ( .A1(n482), .A2(n495), .ZN(n475) );
  NAND2_X1 U524 ( .A1(n475), .A2(n508), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n470), .B(n469), .ZN(G1324GAT) );
  NAND2_X1 U526 ( .A1(n510), .A2(n475), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n471), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U528 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n473) );
  NAND2_X1 U529 ( .A1(n475), .A2(n522), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(G15GAT), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U532 ( .A1(n475), .A2(n524), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  NAND2_X1 U535 ( .A1(n560), .A2(n477), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT101), .B(n478), .Z(n479) );
  NOR2_X1 U537 ( .A1(n578), .A2(n479), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n507) );
  NOR2_X1 U540 ( .A1(n482), .A2(n507), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT104), .B(KEYINPUT38), .Z(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT103), .B(n483), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n492) );
  NAND2_X1 U544 ( .A1(n492), .A2(n508), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(G36GAT), .B(KEYINPUT105), .Z(n489) );
  NAND2_X1 U547 ( .A1(n492), .A2(n510), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n492), .A2(n522), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n524), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U554 ( .A(n565), .ZN(n540) );
  NOR2_X1 U555 ( .A1(n540), .A2(n554), .ZN(n494) );
  XOR2_X1 U556 ( .A(KEYINPUT106), .B(n494), .Z(n506) );
  NOR2_X1 U557 ( .A1(n506), .A2(n495), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT107), .B(n496), .Z(n501) );
  NAND2_X1 U559 ( .A1(n501), .A2(n508), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT42), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n510), .A2(n501), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U564 ( .A1(n501), .A2(n522), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U567 ( .A1(n501), .A2(n524), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT109), .Z(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NOR2_X1 U571 ( .A1(n507), .A2(n506), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n515), .A2(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n510), .A2(n515), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT110), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G92GAT), .B(n512), .ZN(G1337GAT) );
  XOR2_X1 U577 ( .A(G99GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U578 ( .A1(n515), .A2(n522), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n524), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G106GAT), .B(n518), .Z(G1339GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U585 ( .A(n521), .B(KEYINPUT113), .Z(n539) );
  AND2_X1 U586 ( .A1(n522), .A2(n539), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT114), .ZN(n526) );
  INV_X1 U588 ( .A(n524), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n534) );
  NOR2_X1 U590 ( .A1(n565), .A2(n534), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  NOR2_X1 U593 ( .A1(n554), .A2(n534), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  NOR2_X1 U596 ( .A1(n560), .A2(n534), .ZN(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n533), .Z(G1342GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n538), .Z(G1343GAT) );
  NAND2_X1 U604 ( .A1(n563), .A2(n539), .ZN(n549) );
  INV_X1 U605 ( .A(n549), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n540), .A2(n547), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n543) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(n544), .Z(n546) );
  OR2_X1 U612 ( .A1(n549), .A2(n554), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n547), .A2(n573), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U618 ( .A1(n561), .A2(n565), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT121), .ZN(G1348GAT) );
  NOR2_X1 U621 ( .A1(n561), .A2(n554), .ZN(n559) );
  XOR2_X1 U622 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n577), .A2(n565), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U636 ( .A(n577), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

