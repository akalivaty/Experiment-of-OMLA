//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(new_n209), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(new_n218), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n218), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n207), .A2(new_n252), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n249), .B1(new_n250), .B2(new_n251), .C1(new_n201), .C2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(new_n215), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT11), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n248), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT12), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n254), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n261), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n206), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G68), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n260), .A2(new_n264), .A3(new_n265), .A4(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G274), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n230), .A2(G1698), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G226), .B2(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n278), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n277), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G238), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n275), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n291), .B2(new_n290), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n287), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(G169), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n295), .A2(G179), .A3(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n298), .B2(G169), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n270), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(new_n270), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n298), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT73), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n316), .A2(new_n250), .B1(new_n207), .B2(new_n251), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n257), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n268), .A2(G77), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n318), .B1(G77), .B2(new_n261), .C1(new_n266), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G244), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n276), .B1(new_n321), .B2(new_n290), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n281), .A2(new_n283), .A3(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT68), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT3), .B(G33), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT68), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(G1698), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n288), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(G232), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G107), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G107), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n331), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n323), .B1(new_n339), .B2(new_n275), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n320), .B1(new_n340), .B2(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n307), .B2(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n323), .C1(new_n339), .C2(new_n275), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n346), .A3(new_n320), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G223), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n325), .B2(new_n328), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n326), .A2(G222), .A3(new_n330), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n251), .B2(new_n326), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n286), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n290), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n277), .B1(G226), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n313), .A2(new_n250), .B1(new_n359), .B2(new_n253), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT69), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT69), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(new_n359), .B2(new_n253), .C1(new_n313), .C2(new_n250), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n257), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n268), .A2(G50), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n266), .A2(new_n367), .B1(G50), .B2(new_n261), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(KEYINPUT9), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n371));
  INV_X1    g0171(.A(new_n364), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n360), .B2(KEYINPUT69), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n256), .B1(new_n373), .B2(new_n363), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n371), .B1(new_n374), .B2(new_n368), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n354), .A2(G190), .A3(new_n356), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n358), .A2(new_n370), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n368), .B1(new_n365), .B2(new_n257), .ZN(new_n379));
  AOI22_X1  g0179(.A1(G200), .A2(new_n357), .B1(new_n379), .B2(KEYINPUT9), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT10), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(new_n376), .A4(new_n375), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n357), .A2(new_n343), .ZN(new_n384));
  INV_X1    g0184(.A(new_n379), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n354), .A2(new_n345), .A3(new_n356), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n313), .B1(new_n206), .B2(G20), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n267), .A2(new_n390), .B1(new_n313), .B2(new_n262), .ZN(new_n391));
  XNOR2_X1  g0191(.A(G58), .B(G68), .ZN(new_n392));
  INV_X1    g0192(.A(new_n253), .ZN(new_n393));
  AOI22_X1  g0193(.A1(G20), .A2(new_n392), .B1(new_n393), .B2(G159), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT74), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT74), .B1(new_n281), .B2(new_n283), .ZN(new_n396));
  NOR2_X1   g0196(.A1(KEYINPUT7), .A2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n281), .B2(new_n283), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT16), .B(new_n394), .C1(new_n399), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n257), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n281), .A2(new_n283), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n207), .B1(new_n281), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT7), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n400), .A2(new_n401), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(G68), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT16), .B1(new_n410), .B2(new_n394), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n391), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n350), .A2(new_n330), .ZN(new_n413));
  INV_X1    g0213(.A(G226), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G1698), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n281), .A2(new_n413), .A3(new_n283), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n286), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n275), .A2(G232), .A3(new_n289), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n276), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(G169), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n275), .B1(new_n416), .B2(new_n417), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n276), .A2(new_n420), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(G179), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT76), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n421), .A3(new_n345), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n343), .B1(new_n423), .B2(new_n424), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n389), .B1(new_n412), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G200), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n419), .B2(new_n421), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT77), .B(G190), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n423), .A2(new_n424), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n391), .C1(new_n404), .C2(new_n411), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n412), .A2(new_n431), .A3(new_n389), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n440), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n433), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n349), .A2(new_n388), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n310), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT25), .B1(new_n262), .B2(new_n332), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n332), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n206), .A2(G33), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n261), .A2(new_n450), .A3(new_n215), .A4(new_n255), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n448), .A2(new_n449), .B1(G107), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n326), .A2(G257), .A3(G1698), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G294), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n326), .A2(G250), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(G1698), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n286), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n272), .A2(G1), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(G274), .A3(new_n275), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n286), .B1(new_n460), .B2(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G264), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n434), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n457), .A2(new_n286), .B1(G264), .B2(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n307), .A3(new_n461), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n281), .A2(new_n283), .A3(new_n207), .A4(G87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT22), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n326), .A2(new_n471), .A3(new_n207), .A4(G87), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n332), .A3(G20), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n474), .A2(new_n332), .A3(KEYINPUT85), .A4(G20), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n333), .A2(new_n335), .A3(G20), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT80), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G116), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n207), .A3(G33), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT24), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n470), .A2(new_n472), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n252), .B1(new_n484), .B2(new_n486), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n207), .A2(new_n492), .B1(new_n480), .B2(new_n481), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n479), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT86), .B1(new_n496), .B2(new_n257), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT86), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n498), .B(new_n256), .C1(new_n490), .C2(new_n495), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n453), .B(new_n468), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n453), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n498), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(KEYINPUT86), .A3(new_n257), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n464), .A2(G179), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n343), .B2(new_n464), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n500), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n451), .A2(new_n483), .B1(new_n261), .B2(new_n487), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n485), .A2(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n483), .A2(KEYINPUT80), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n256), .B1(new_n514), .B2(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n207), .C1(G33), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n252), .A2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n207), .A4(new_n516), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n515), .A2(new_n523), .A3(KEYINPUT20), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT20), .B1(new_n515), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n511), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n459), .A2(new_n460), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(G270), .A3(new_n275), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n529), .A2(new_n461), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n326), .A2(G257), .A3(new_n330), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n326), .A2(G264), .A3(G1698), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n284), .A2(G303), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n286), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n527), .A2(KEYINPUT21), .A3(G169), .A4(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(G169), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n515), .A2(new_n523), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n510), .B1(new_n542), .B2(new_n524), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n538), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n530), .A2(new_n535), .A3(G179), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n527), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n536), .A2(G200), .ZN(new_n547));
  INV_X1    g0347(.A(new_n436), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n530), .A2(new_n535), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  AND4_X1   g0350(.A1(new_n537), .A2(new_n544), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n261), .A2(G97), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n452), .B2(G97), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n408), .A2(new_n409), .A3(new_n336), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n517), .A2(new_n332), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n332), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G20), .B1(G77), .B2(new_n393), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT78), .B1(new_n562), .B2(new_n257), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT78), .ZN(new_n564));
  AOI211_X1 g0364(.A(new_n564), .B(new_n256), .C1(new_n554), .C2(new_n561), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n553), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(new_n281), .A3(new_n283), .A4(G244), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n516), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT4), .B1(new_n326), .B2(G244), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G250), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n284), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(G1698), .B1(new_n575), .B2(new_n568), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n275), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n528), .A2(G257), .A3(new_n275), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n345), .A3(new_n461), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n567), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n568), .B1(new_n284), .B2(new_n321), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n516), .A3(new_n570), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n330), .B1(new_n456), .B2(KEYINPUT4), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n286), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n578), .A2(new_n461), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(KEYINPUT79), .A3(new_n345), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n580), .A2(new_n586), .B1(new_n343), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n566), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n562), .A2(new_n257), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n564), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n562), .A2(KEYINPUT78), .A3(new_n257), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n584), .A2(G190), .A3(new_n585), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n434), .B1(new_n584), .B2(new_n585), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n596), .A3(new_n553), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G87), .A2(G97), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n333), .A2(new_n335), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n207), .B1(new_n278), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n600), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n281), .A2(new_n283), .A3(new_n207), .A4(G68), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n602), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n257), .ZN(new_n610));
  INV_X1    g0410(.A(new_n316), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n261), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n452), .A2(G87), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G33), .B1(new_n512), .B2(new_n513), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n288), .A2(new_n330), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n321), .A2(G1698), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n281), .A2(new_n617), .A3(new_n283), .A4(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n275), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G274), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n460), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n574), .B1(new_n272), .B2(G1), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n275), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(G200), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(G238), .A2(G1698), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n321), .B2(G1698), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n326), .B1(new_n487), .B2(G33), .ZN(new_n629));
  OAI211_X1 g0429(.A(G190), .B(new_n624), .C1(new_n629), .C2(new_n275), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n615), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n612), .B1(new_n609), .B2(new_n257), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT82), .B1(new_n452), .B2(new_n611), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT82), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n451), .A2(new_n635), .A3(new_n316), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(G169), .B1(new_n620), .B2(new_n625), .ZN(new_n638));
  OAI211_X1 g0438(.A(G179), .B(new_n624), .C1(new_n629), .C2(new_n275), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n633), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n551), .A2(new_n589), .A3(new_n597), .A4(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n446), .A2(new_n509), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n387), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n412), .A2(new_n431), .A3(new_n389), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n432), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n347), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n347), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n308), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n304), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n439), .B(KEYINPUT17), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n654), .A2(new_n655), .B1(new_n378), .B2(new_n382), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n644), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n632), .A2(new_n640), .A3(KEYINPUT87), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT87), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n633), .A2(new_n637), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n638), .A2(new_n639), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n633), .A2(new_n614), .A3(new_n626), .A4(new_n630), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n500), .A3(new_n589), .A4(new_n597), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n544), .A2(new_n537), .A3(new_n546), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n453), .B1(new_n497), .B2(new_n499), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n507), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n566), .A2(new_n641), .A3(new_n588), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT87), .B1(new_n632), .B2(new_n640), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n663), .A2(new_n660), .A3(new_n664), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n566), .A3(new_n588), .A4(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n673), .B(new_n663), .C1(KEYINPUT26), .C2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n658), .B1(new_n446), .B2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT90), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT27), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT90), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n206), .A3(new_n207), .A4(G13), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT91), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n681), .A2(KEYINPUT91), .A3(new_n682), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G213), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n684), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n543), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n668), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n544), .A2(new_n537), .A3(new_n550), .A4(new_n546), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n505), .A2(new_n696), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n669), .A2(new_n507), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n509), .A2(new_n702), .B1(new_n703), .B2(new_n696), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n703), .A2(new_n500), .ZN(new_n706));
  INV_X1    g0506(.A(new_n668), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n695), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n669), .A2(new_n507), .A3(new_n696), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n705), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n210), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G1), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n337), .A2(new_n483), .A3(new_n598), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(new_n213), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n597), .A2(new_n589), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n699), .A2(new_n640), .A3(new_n632), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n706), .A2(new_n721), .A3(new_n722), .A4(new_n696), .ZN(new_n723));
  INV_X1    g0523(.A(new_n587), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n620), .A2(new_n625), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n458), .A2(new_n463), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n724), .A2(new_n726), .A3(new_n545), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n725), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n587), .A2(new_n464), .A3(new_n536), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n466), .A2(new_n725), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n530), .A2(new_n535), .A3(G179), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n729), .B1(new_n736), .B2(new_n724), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n695), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT31), .B(new_n695), .C1(new_n733), .C2(new_n737), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n720), .B1(new_n723), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n696), .B1(new_n671), .B2(new_n677), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT93), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT93), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n696), .C1(new_n671), .C2(new_n677), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT26), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n566), .A2(new_n641), .A3(new_n588), .A4(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n750), .A2(new_n663), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n703), .A2(new_n707), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n674), .A2(new_n675), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n505), .B2(new_n468), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n756), .A3(new_n721), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n695), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT29), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n743), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n719), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(G13), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G45), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n716), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n215), .B1(G20), .B2(new_n343), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n207), .B1(new_n774), .B2(G190), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n775), .A2(KEYINPUT100), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(KEYINPUT100), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n517), .ZN(new_n780));
  NAND2_X1  g0580(.A1(G20), .A2(G179), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n434), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n436), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n548), .A3(G200), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n202), .B1(new_n201), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n783), .A2(G190), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n780), .B(new_n787), .C1(G77), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n345), .A2(G200), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n307), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n332), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n207), .A2(new_n307), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n284), .B(new_n795), .C1(G87), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n793), .A2(new_n774), .ZN(new_n800));
  INV_X1    g0600(.A(G159), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n782), .A2(new_n307), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT99), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G68), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n789), .A2(new_n799), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n779), .A2(new_n812), .B1(new_n785), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n788), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  INV_X1    g0616(.A(G326), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n815), .A2(new_n816), .B1(new_n817), .B2(new_n786), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT33), .B(G317), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n809), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n797), .B(KEYINPUT101), .Z(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G303), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n284), .B1(new_n794), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n800), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G329), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n819), .A2(new_n821), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n773), .B1(new_n811), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G13), .A2(G33), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(G20), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n772), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n395), .A2(new_n396), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n713), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n272), .B2(new_n214), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n243), .B2(new_n272), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n713), .A2(new_n284), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(G355), .B1(new_n483), .B2(new_n713), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n771), .B(new_n829), .C1(new_n833), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n832), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n700), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT102), .ZN(new_n846));
  INV_X1    g0646(.A(new_n771), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n701), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(G330), .B2(new_n700), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(G396));
  NAND4_X1  g0650(.A1(new_n649), .A2(new_n320), .A3(new_n650), .A4(new_n695), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n320), .A2(new_n695), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n342), .A2(new_n347), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n745), .A2(new_n748), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n854), .B(new_n696), .C1(new_n671), .C2(new_n677), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n743), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n769), .B2(new_n770), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(new_n743), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n772), .A2(new_n830), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n847), .B1(G77), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n786), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G143), .A2(new_n784), .B1(new_n865), .B2(G137), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n866), .B1(new_n801), .B2(new_n815), .C1(new_n808), .C2(new_n359), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT34), .Z(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n835), .B1(new_n800), .B2(new_n869), .C1(new_n248), .C2(new_n794), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(G58), .B2(new_n778), .ZN(new_n871));
  INV_X1    g0671(.A(new_n822), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n201), .B2(new_n872), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n812), .A2(new_n785), .B1(new_n815), .B2(new_n514), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n780), .B(new_n874), .C1(G303), .C2(new_n865), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n284), .B1(new_n800), .B2(new_n816), .ZN(new_n876));
  INV_X1    g0676(.A(new_n794), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(G87), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n875), .B(new_n878), .C1(new_n332), .C2(new_n872), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n808), .A2(new_n824), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n868), .A2(new_n873), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n864), .B1(new_n881), .B2(new_n772), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n831), .B2(new_n854), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n861), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  OR2_X1    g0685(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n216), .A4(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(G77), .B1(new_n202), .B2(new_n248), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n892), .A2(new_n213), .B1(G50), .B2(new_n248), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(G1), .A3(new_n762), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT104), .ZN(new_n896));
  INV_X1    g0696(.A(new_n446), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n749), .A2(new_n897), .A3(new_n759), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n658), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n412), .A2(new_n431), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT107), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n689), .A2(new_n903), .A3(new_n692), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n689), .B2(new_n692), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n412), .A2(new_n906), .ZN(new_n907));
  AND4_X1   g0707(.A1(new_n901), .A2(new_n902), .A3(new_n907), .A4(new_n439), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n284), .A2(new_n207), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n248), .B1(new_n909), .B2(KEYINPUT7), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT74), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n284), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n326), .A2(KEYINPUT74), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(new_n397), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT16), .B1(new_n915), .B2(new_n394), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n391), .B1(new_n404), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n693), .ZN(new_n920));
  OAI211_X1 g0720(.A(KEYINPUT106), .B(new_n391), .C1(new_n404), .C2(new_n916), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(new_n431), .A3(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n439), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n908), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n922), .B1(new_n646), .B2(new_n653), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n444), .A2(new_n412), .A3(new_n906), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n902), .A2(new_n907), .A3(new_n439), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT37), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n902), .A2(new_n907), .A3(new_n901), .A4(new_n439), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT38), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n900), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n927), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(KEYINPUT38), .C1(new_n937), .C2(new_n908), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n926), .B1(new_n925), .B2(new_n927), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(KEYINPUT39), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n302), .A2(new_n303), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n270), .A3(new_n696), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n935), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n695), .A2(new_n270), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n304), .A2(new_n308), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n270), .B(new_n695), .C1(new_n302), .C2(new_n303), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n347), .A2(new_n695), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n857), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n938), .A2(new_n939), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n646), .A2(new_n906), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n944), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n899), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n740), .A2(new_n741), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n642), .A2(new_n509), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(new_n696), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n949), .A2(new_n854), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT108), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n723), .A2(new_n742), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n947), .A2(new_n948), .B1(new_n851), .B2(new_n853), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT40), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT108), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n963), .A2(new_n968), .A3(new_n954), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n928), .A2(new_n934), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n642), .A2(new_n509), .A3(new_n695), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n965), .B1(new_n971), .B2(new_n959), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT40), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n446), .A2(new_n961), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n720), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n958), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n206), .B2(new_n763), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n958), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n896), .B1(new_n979), .B2(new_n980), .ZN(G367));
  INV_X1    g0781(.A(KEYINPUT113), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n566), .A2(new_n695), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n721), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n566), .A2(new_n588), .A3(new_n695), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n705), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT110), .Z(new_n988));
  INV_X1    g0788(.A(KEYINPUT112), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n706), .A3(new_n708), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT109), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n589), .B1(new_n984), .B2(new_n703), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n991), .A2(KEYINPUT42), .B1(new_n696), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n695), .A2(new_n615), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n666), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n663), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n993), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n990), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n998), .B(KEYINPUT43), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n993), .B2(new_n995), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT111), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n988), .A2(new_n989), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n988), .A2(new_n989), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n766), .A2(new_n206), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n986), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n711), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT44), .Z(new_n1016));
  NOR2_X1   g0816(.A1(new_n711), .A2(new_n1014), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(new_n705), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(new_n701), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n760), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n714), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1013), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n982), .B1(new_n1011), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n760), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n705), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1019), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1022), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1012), .B1(new_n1032), .B2(new_n1024), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1033), .A2(KEYINPUT113), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n833), .B1(new_n210), .B2(new_n316), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n836), .B2(new_n236), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n771), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n815), .A2(new_n201), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n779), .A2(new_n248), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G143), .C2(new_n865), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G58), .A2(new_n798), .B1(new_n826), .B2(G137), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT114), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n877), .A2(G77), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n326), .C1(new_n359), .C2(new_n785), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n809), .A2(G159), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1041), .A2(new_n1044), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n877), .A2(G97), .ZN(new_n1050));
  INV_X1    g0850(.A(G317), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n834), .C1(new_n1051), .C2(new_n800), .ZN(new_n1052));
  INV_X1    g0852(.A(G303), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n824), .A2(new_n815), .B1(new_n785), .B2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n779), .A2(new_n337), .B1(new_n786), .B2(new_n816), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n812), .B2(new_n808), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n514), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n822), .A2(G116), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(KEYINPUT46), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT47), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n1038), .B1(new_n844), .B2(new_n998), .C1(new_n1062), .C2(new_n773), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1035), .A2(new_n1063), .ZN(G387));
  OR2_X1    g0864(.A1(new_n704), .A2(new_n844), .ZN(new_n1065));
  AOI211_X1 g0865(.A(G45), .B(new_n717), .C1(G68), .C2(G77), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n313), .A2(G50), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT50), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n837), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n272), .B2(new_n233), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n840), .A2(new_n717), .B1(new_n332), .B2(new_n713), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT115), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n833), .B1(new_n1072), .B2(KEYINPUT115), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n847), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1050), .B(new_n835), .C1(new_n248), .C2(new_n815), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n251), .A2(new_n797), .B1(new_n800), .B2(new_n359), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1077), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n778), .A2(new_n611), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n801), .B2(new_n786), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G50), .B2(new_n784), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n313), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n809), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n779), .A2(new_n824), .B1(new_n812), .B2(new_n797), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n788), .A2(G303), .B1(new_n865), .B2(G322), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n1051), .B2(new_n785), .C1(new_n808), .C2(new_n816), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT49), .Z(new_n1093));
  OAI221_X1 g0893(.A(new_n834), .B1(new_n800), .B2(new_n817), .C1(new_n514), .C2(new_n794), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1086), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1075), .B1(new_n1095), .B2(new_n772), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1031), .A2(new_n1013), .B1(new_n1065), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1031), .A2(new_n760), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n714), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1031), .A2(new_n760), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(G393));
  AND2_X1   g0901(.A1(new_n1020), .A2(new_n1098), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n714), .B1(new_n1020), .B2(new_n1098), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1014), .A2(new_n832), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n833), .B1(new_n517), .B2(new_n210), .C1(new_n837), .C2(new_n246), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n847), .A2(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n785), .A2(new_n816), .B1(new_n1051), .B2(new_n786), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT52), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n779), .A2(new_n514), .B1(new_n815), .B2(new_n812), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n824), .A2(new_n797), .B1(new_n800), .B2(new_n813), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n1110), .A2(new_n326), .A3(new_n795), .A4(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1112), .C1(new_n1053), .C2(new_n808), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G68), .A2(new_n798), .B1(new_n826), .B2(G143), .ZN(new_n1114));
  INV_X1    g0914(.A(G87), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1114), .B(new_n835), .C1(new_n1115), .C2(new_n794), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT117), .Z(new_n1117));
  OAI22_X1  g0917(.A1(new_n785), .A2(new_n801), .B1(new_n359), .B2(new_n786), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n778), .A2(G77), .B1(new_n788), .B2(new_n1084), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n201), .C2(new_n808), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1113), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1107), .B1(new_n1122), .B2(new_n772), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1030), .A2(new_n1013), .B1(new_n1105), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1104), .A2(new_n1124), .ZN(G390));
  NAND2_X1  g0925(.A1(new_n897), .A2(new_n743), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n898), .A2(new_n658), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n854), .C1(new_n971), .C2(new_n959), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n950), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n964), .A2(G330), .A3(new_n854), .A4(new_n949), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n951), .B1(new_n758), .B2(new_n854), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n663), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n673), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n695), .B1(new_n1137), .B2(new_n757), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n951), .B1(new_n1138), .B2(new_n854), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1128), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n750), .A2(new_n663), .A3(new_n752), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n854), .B(new_n696), .C1(new_n671), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n952), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n949), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n929), .A2(new_n933), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n926), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n943), .B1(new_n1148), .B2(new_n938), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n950), .B1(new_n1143), .B2(new_n952), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n942), .B1(new_n928), .B2(new_n934), .ZN(new_n1152));
  OAI21_X1  g0952(.A(KEYINPUT118), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n935), .A2(new_n940), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n943), .B2(new_n953), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1154), .A2(new_n1156), .A3(new_n1131), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1131), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1141), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1141), .B(KEYINPUT119), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1146), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT118), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1156), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1129), .A2(new_n950), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1154), .A2(new_n1156), .A3(new_n1131), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1139), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(new_n1127), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1161), .A2(new_n714), .A3(new_n1162), .A4(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n788), .A2(new_n1176), .B1(new_n784), .B2(G132), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n284), .B1(new_n826), .B2(G125), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n201), .C2(new_n794), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n797), .A2(new_n359), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n786), .C1(new_n801), .C2(new_n779), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1179), .B(new_n1184), .C1(G137), .C2(new_n809), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n284), .B1(new_n251), .B2(new_n779), .C1(new_n872), .C2(new_n1115), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n794), .A2(new_n248), .B1(new_n800), .B2(new_n812), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT121), .Z(new_n1188));
  AOI22_X1  g0988(.A1(G116), .A2(new_n784), .B1(new_n865), .B2(G283), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n517), .B2(new_n815), .C1(new_n808), .C2(new_n337), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n772), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n847), .C1(new_n1084), .C2(new_n863), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1155), .B2(new_n830), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n1013), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1174), .A2(new_n1196), .ZN(G378));
  INV_X1    g0997(.A(new_n957), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n379), .A2(new_n693), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n388), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1199), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n383), .A2(new_n387), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1203), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1201), .B1(new_n383), .B2(new_n387), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1199), .B(new_n644), .C1(new_n378), .C2(new_n382), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1204), .A2(new_n1208), .A3(KEYINPUT123), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT123), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n720), .B(new_n1211), .C1(new_n973), .C2(new_n969), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n974), .B2(G330), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1198), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1211), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n974), .A2(G330), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n720), .B1(new_n969), .B2(new_n973), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n957), .C1(new_n1219), .C2(new_n1214), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1173), .A2(new_n1128), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n715), .B1(new_n1221), .B2(KEYINPUT57), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1127), .B1(new_n1195), .B2(new_n1172), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n332), .A2(new_n785), .B1(new_n815), .B2(new_n316), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1040), .B(new_n1228), .C1(G116), .C2(new_n865), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n834), .A2(new_n271), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n794), .A2(new_n202), .B1(new_n800), .B2(new_n824), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(G77), .C2(new_n798), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1229), .B(new_n1232), .C1(new_n517), .C2(new_n808), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT58), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1230), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G137), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n815), .A2(new_n1239), .B1(new_n797), .B2(new_n1175), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n778), .A2(G150), .B1(new_n865), .B2(G125), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1183), .B2(new_n785), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G132), .C2(new_n809), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT59), .Z(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(KEYINPUT122), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n826), .C2(G124), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n801), .B2(new_n794), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1244), .B2(KEYINPUT122), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1235), .B(new_n1238), .C1(new_n1245), .C2(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n847), .B1(G50), .B2(new_n863), .C1(new_n1249), .C2(new_n773), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n830), .B2(new_n1217), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1013), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1227), .A2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n1171), .A2(new_n1127), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1141), .A2(new_n1025), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1140), .A2(new_n1013), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n771), .B1(new_n248), .B2(new_n862), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n822), .A2(G159), .B1(G128), .B2(new_n826), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT124), .Z(new_n1260));
  OAI221_X1 g1060(.A(new_n835), .B1(new_n202), .B2(new_n794), .C1(new_n815), .C2(new_n359), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n778), .A2(G50), .B1(new_n865), .B2(G132), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1239), .B2(new_n785), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(new_n809), .C2(new_n1176), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n809), .A2(new_n487), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1045), .B(new_n284), .C1(new_n1053), .C2(new_n800), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n788), .A2(new_n336), .B1(new_n784), .B2(G283), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1267), .B(new_n1081), .C1(new_n812), .C2(new_n786), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(G97), .C2(new_n822), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1260), .A2(new_n1264), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1258), .B1(new_n1270), .B2(new_n773), .C1(new_n949), .C2(new_n831), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1257), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1256), .A2(new_n1273), .ZN(G381));
  INV_X1    g1074(.A(G390), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1035), .A2(new_n1063), .A3(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1276), .A2(G384), .A3(G381), .A4(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1174), .A2(KEYINPUT125), .A3(new_n1196), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT125), .B1(new_n1174), .B2(new_n1196), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1253), .A3(new_n1227), .A4(new_n1281), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n694), .A2(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(G375), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1281), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(G213), .A3(new_n1285), .ZN(G409));
  XOR2_X1   g1086(.A(G393), .B(G396), .Z(new_n1287));
  AND3_X1   g1087(.A1(new_n1035), .A2(new_n1063), .A3(new_n1275), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1275), .B1(new_n1035), .B2(new_n1063), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(G390), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1287), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1276), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT60), .B1(new_n1171), .B2(new_n1127), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n715), .B1(new_n1295), .B2(new_n1255), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1171), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1296), .A2(KEYINPUT126), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT126), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1273), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n884), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G384), .B(new_n1273), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1173), .A2(new_n1128), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1025), .A3(new_n1252), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1253), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1279), .A2(new_n1280), .A3(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1227), .A2(G378), .A3(new_n1253), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1283), .B(new_n1303), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1280), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1174), .A2(KEYINPUT125), .A3(new_n1196), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1306), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1227), .A2(G378), .A3(new_n1253), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1317), .A2(KEYINPUT62), .A3(new_n1283), .A4(new_n1303), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1312), .A2(KEYINPUT127), .A3(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1283), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n694), .A2(G213), .A3(G2897), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1301), .A2(new_n1302), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1310), .A2(new_n1326), .A3(new_n1311), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1294), .B1(new_n1319), .B2(new_n1328), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1310), .A2(new_n1331), .ZN(new_n1332));
  OR2_X1    g1132(.A1(new_n1310), .A2(new_n1331), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1330), .A2(new_n1325), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1329), .A2(new_n1334), .ZN(G405));
  AOI21_X1  g1135(.A(new_n1309), .B1(G375), .B2(new_n1281), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1303), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1330), .B(new_n1337), .ZN(G402));
endmodule


