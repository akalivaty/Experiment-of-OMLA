//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT10), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(KEYINPUT65), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n191), .A2(KEYINPUT65), .A3(G146), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n191), .B2(G146), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n199), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n197), .A2(KEYINPUT67), .A3(new_n202), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n201), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n190), .B1(new_n209), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n223));
  INV_X1    g037(.A(G134), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G137), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT11), .A3(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n225), .A3(new_n227), .A4(new_n228), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n191), .A2(G146), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n199), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n200), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n195), .A2(new_n196), .ZN(new_n241));
  AND4_X1   g055(.A1(KEYINPUT67), .A2(new_n241), .A3(new_n199), .A4(new_n202), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n197), .B2(new_n202), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n221), .A2(new_n190), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT78), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT4), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n215), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n247), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT0), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(new_n198), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n199), .A2(new_n237), .B1(KEYINPUT0), .B2(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n198), .A3(KEYINPUT64), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(KEYINPUT0), .B2(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n197), .A2(new_n259), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n247), .A2(G101), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n257), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n222), .A2(new_n236), .A3(new_n246), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n197), .A2(new_n200), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n242), .B2(new_n243), .ZN(new_n272));
  INV_X1    g086(.A(new_n221), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n240), .B(new_n221), .C1(new_n242), .C2(new_n243), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n270), .B(new_n236), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n209), .B2(new_n221), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT12), .B1(new_n277), .B2(new_n235), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n269), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n269), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n257), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n267), .A2(new_n265), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n239), .B1(new_n207), .B2(new_n208), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(KEYINPUT10), .ZN(new_n289));
  OAI22_X1  g103(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT10), .B1(new_n272), .B2(new_n273), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n235), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n279), .A2(new_n283), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G469), .B1(new_n293), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n276), .A2(new_n278), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n269), .A2(new_n284), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n284), .B1(new_n292), .B2(new_n269), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n295), .B(new_n296), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G113), .B(G122), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(new_n210), .ZN(new_n304));
  OR2_X1    g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(G143), .A2(G214), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n230), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  AOI21_X1  g122(.A(G143), .B1(new_n308), .B2(G214), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT89), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G214), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n191), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n230), .A4(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n305), .A2(new_n306), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n316), .B2(new_n309), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n322), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT19), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n318), .B(new_n325), .C1(G146), .C2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n194), .B1(new_n320), .B2(new_n322), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n322), .A3(new_n194), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT88), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n320), .A2(new_n322), .A3(new_n194), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n312), .A2(KEYINPUT18), .A3(G131), .A4(new_n314), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT18), .A2(G131), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n316), .B2(new_n309), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n304), .B1(new_n328), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n310), .A2(new_n315), .A3(new_n317), .A4(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n323), .A2(new_n324), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n194), .ZN(new_n348));
  OAI211_X1 g162(.A(KEYINPUT17), .B(G131), .C1(new_n316), .C2(new_n309), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n325), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n341), .B(new_n304), .C1(new_n346), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n348), .A2(new_n325), .A3(new_n349), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n354), .A2(new_n345), .B1(new_n336), .B2(new_n340), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT90), .B1(new_n355), .B2(new_n304), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n343), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n352), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(KEYINPUT90), .A3(new_n304), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n342), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT92), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT91), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(KEYINPUT91), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n359), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(KEYINPUT20), .B2(new_n372), .ZN(new_n373));
  OAI22_X1  g187(.A1(new_n353), .A2(new_n356), .B1(new_n304), .B2(new_n355), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n296), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n375), .A2(G475), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT93), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n378));
  INV_X1    g192(.A(new_n376), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n366), .A2(KEYINPUT91), .ZN(new_n380));
  AOI211_X1 g194(.A(new_n369), .B(new_n342), .C1(new_n364), .C2(new_n365), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n360), .B1(new_n382), .B2(new_n359), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n378), .B(new_n379), .C1(new_n383), .C2(new_n368), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n191), .A2(G128), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n198), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n224), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT94), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G116), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n213), .B1(new_n393), .B2(KEYINPUT14), .ZN(new_n394));
  XNOR2_X1  g208(.A(G116), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n397), .A3(new_n389), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n385), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n386), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n385), .A2(new_n400), .ZN(new_n403));
  OAI21_X1  g217(.A(G134), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n395), .A2(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(G107), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n389), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n187), .A2(new_n408), .A3(G953), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n399), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n399), .B2(new_n407), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n296), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G478), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(KEYINPUT15), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT95), .B(new_n296), .C1(new_n410), .C2(new_n411), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n412), .A2(new_n416), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G952), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n421), .A2(KEYINPUT96), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(KEYINPUT96), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n281), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(G234), .A2(G237), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G898), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n281), .B1(KEYINPUT21), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(KEYINPUT21), .B2(new_n428), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(G902), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n420), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n377), .A2(new_n384), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT87), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G113), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G116), .B(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT5), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT2), .B(G113), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n443), .A2(new_n445), .B1(new_n447), .B2(new_n444), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n273), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n444), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n440), .A2(G116), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n446), .B1(new_n441), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n256), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n255), .B1(new_n247), .B2(new_n252), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n267), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n449), .B1(new_n456), .B2(KEYINPUT80), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n459), .A2(new_n266), .B1(new_n450), .B2(new_n452), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n460), .B2(new_n257), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n438), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n458), .A3(new_n257), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n437), .A4(new_n449), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(KEYINPUT6), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n288), .A2(new_n321), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n265), .A2(new_n321), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G224), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT82), .B1(new_n470), .B2(G953), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n281), .A3(G224), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT81), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT83), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n469), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n438), .C1(new_n457), .C2(new_n461), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n466), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT7), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n467), .A2(new_n468), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT85), .B(KEYINPUT7), .Z(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n474), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n467), .B2(new_n468), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n217), .A2(new_n220), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n448), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n448), .A2(new_n487), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n437), .B(KEYINPUT8), .Z(new_n490));
  NOR3_X1   g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n482), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n492), .B2(new_n465), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n480), .A2(KEYINPUT86), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT86), .B1(new_n480), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n436), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n493), .A3(new_n435), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n434), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n504));
  INV_X1    g318(.A(new_n453), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n265), .A2(new_n235), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n229), .A2(new_n230), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n226), .A2(G134), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n228), .A3(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT68), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n505), .B(new_n506), .C1(new_n514), .C2(new_n288), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n308), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n265), .A2(new_n235), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n507), .A2(new_n512), .A3(new_n509), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n512), .B1(new_n507), .B2(new_n509), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n525), .B1(new_n528), .B2(new_n244), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n505), .ZN(new_n530));
  INV_X1    g344(.A(new_n515), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT28), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n510), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n506), .B1(new_n288), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n453), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n515), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT70), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n541), .B(new_n538), .C1(new_n536), .C2(new_n515), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n540), .A2(new_n542), .A3(new_n522), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n506), .C1(new_n288), .C2(new_n534), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n529), .B2(new_n544), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n531), .B1(new_n546), .B2(new_n453), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n523), .B1(new_n547), .B2(new_n521), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n533), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G472), .ZN(new_n550));
  NOR2_X1   g364(.A1(G472), .A2(G902), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT32), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n540), .A2(new_n542), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n521), .B1(new_n554), .B2(new_n517), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n244), .A2(new_n511), .A3(new_n513), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n544), .B1(new_n556), .B2(new_n506), .ZN(new_n557));
  INV_X1    g371(.A(new_n545), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n453), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n515), .A3(new_n521), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n547), .A2(new_n562), .A3(new_n521), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n553), .B1(new_n555), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n550), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n517), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n540), .A2(new_n542), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n561), .B(new_n563), .C1(new_n568), .C2(new_n521), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT32), .B1(new_n569), .B2(new_n551), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n504), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n569), .A2(new_n553), .B1(new_n549), .B2(G472), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n551), .B1(new_n555), .B2(new_n564), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT32), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n575), .A3(KEYINPUT71), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G234), .ZN(new_n578));
  OAI21_X1  g392(.A(G217), .B1(new_n578), .B2(G902), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n440), .A2(G128), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n198), .A2(G119), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT24), .B(G110), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT73), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT23), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n440), .B2(G128), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n583), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n588), .B(new_n590), .C1(G110), .C2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n325), .A3(new_n331), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n348), .A2(new_n325), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT72), .A4(new_n583), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(G110), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n597), .B(new_n601), .C1(new_n585), .C2(new_n586), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n596), .A2(new_n602), .A3(KEYINPUT74), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT74), .B1(new_n596), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n582), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n582), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n596), .A2(new_n602), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT74), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT75), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT25), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n605), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n611), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n579), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n614), .B2(new_n613), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n605), .A2(new_n609), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n578), .B2(G217), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT76), .B1(new_n577), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT76), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n623), .B(new_n620), .C1(new_n571), .C2(new_n576), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n302), .B(new_n503), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n569), .B2(new_n296), .ZN(new_n628));
  INV_X1    g442(.A(new_n573), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n621), .A3(new_n302), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n410), .A2(new_n411), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT33), .Z(new_n634));
  NOR2_X1   g448(.A1(new_n415), .A2(G902), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n414), .A2(new_n417), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n634), .A2(new_n635), .B1(new_n636), .B2(new_n415), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n432), .A2(new_n427), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n435), .B1(new_n480), .B2(new_n493), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n501), .B(new_n638), .C1(new_n499), .C2(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n637), .B(new_n640), .C1(new_n377), .C2(new_n384), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n638), .B(KEYINPUT97), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n380), .A2(new_n381), .A3(new_n361), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n379), .B(new_n646), .C1(new_n383), .C2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n501), .B(new_n420), .C1(new_n499), .C2(new_n639), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n420), .A2(new_n501), .ZN(new_n651));
  INV_X1    g465(.A(new_n639), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n498), .ZN(new_n653));
  INV_X1    g467(.A(new_n647), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n372), .A2(KEYINPUT20), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n376), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n653), .A2(new_n656), .A3(KEYINPUT98), .A4(new_n646), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n632), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT99), .Z(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n606), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n607), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n618), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n616), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n630), .A2(new_n302), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n503), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT37), .B(G110), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT100), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(G12));
  AOI21_X1  g485(.A(new_n502), .B1(new_n652), .B2(new_n498), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n672), .A2(new_n302), .A3(new_n666), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n431), .A2(G900), .A3(new_n281), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n427), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n656), .A2(new_n420), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n577), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  INV_X1    g495(.A(KEYINPUT38), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n500), .B(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n521), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n547), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n530), .A2(new_n531), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n627), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n569), .B2(new_n553), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n575), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n651), .A3(new_n666), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n377), .A2(new_n384), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n678), .B(KEYINPUT39), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n302), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT40), .Z(new_n697));
  NAND4_X1  g511(.A1(new_n683), .A2(new_n693), .A3(new_n694), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  INV_X1    g513(.A(new_n678), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n637), .B(new_n700), .C1(new_n377), .C2(new_n384), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n577), .A2(new_n701), .A3(new_n673), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  OR2_X1    g517(.A1(new_n276), .A2(new_n278), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n300), .B1(new_n704), .B2(new_n285), .ZN(new_n705));
  OAI21_X1  g519(.A(G469), .B1(new_n705), .B2(G902), .ZN(new_n706));
  INV_X1    g520(.A(new_n189), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n301), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n577), .A2(new_n641), .A3(new_n621), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n577), .A2(new_n658), .A3(new_n621), .A4(new_n708), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n672), .A3(new_n666), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n434), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n577), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  AND2_X1   g531(.A1(new_n532), .A2(new_n517), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n561), .B(new_n563), .C1(new_n718), .C2(new_n521), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n551), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n706), .A2(new_n707), .A3(new_n301), .A4(new_n646), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n628), .A2(new_n721), .A3(new_n722), .A4(new_n620), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n649), .B1(new_n377), .B2(new_n384), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR2_X1   g540(.A1(new_n628), .A2(new_n721), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n666), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n708), .A2(new_n672), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n701), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n565), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n569), .A2(KEYINPUT103), .A3(new_n553), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n575), .A2(new_n736), .A3(new_n550), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n499), .A2(new_n502), .ZN(new_n739));
  AND4_X1   g553(.A1(KEYINPUT42), .A2(new_n302), .A3(new_n496), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n621), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n637), .B1(new_n377), .B2(new_n384), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n678), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n734), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n562), .B1(new_n547), .B2(new_n521), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n537), .A2(new_n539), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n541), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n537), .A2(KEYINPUT70), .A3(new_n539), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n517), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n684), .ZN(new_n752));
  AOI211_X1 g566(.A(new_n735), .B(new_n552), .C1(new_n747), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT103), .B1(new_n569), .B2(new_n553), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n573), .A2(new_n574), .B1(G472), .B2(new_n549), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n620), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n701), .A3(KEYINPUT104), .A4(new_n740), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n496), .A2(new_n739), .ZN(new_n759));
  INV_X1    g573(.A(new_n302), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n760), .A3(new_n620), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n577), .A2(new_n701), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n763));
  AOI22_X1  g577(.A1(new_n744), .A2(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(KEYINPUT105), .B(G131), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G33));
  NOR3_X1   g580(.A1(new_n566), .A2(new_n570), .A3(new_n504), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT71), .B1(new_n572), .B2(new_n575), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n761), .B(new_n679), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n637), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n377), .A2(new_n384), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n630), .A2(new_n729), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(KEYINPUT44), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT106), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT44), .B1(new_n776), .B2(new_n777), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n293), .A2(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n293), .B2(KEYINPUT45), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(G469), .A2(G902), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n784), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n301), .A3(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n789), .A2(new_n707), .A3(new_n695), .ZN(new_n790));
  INV_X1    g604(.A(new_n759), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n780), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n779), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  NAND2_X1  g609(.A1(new_n789), .A2(new_n707), .ZN(new_n796));
  XOR2_X1   g610(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n791), .A2(new_n620), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n800), .A2(new_n577), .A3(new_n743), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n319), .ZN(G42));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n804));
  NOR2_X1   g618(.A1(G952), .A2(G953), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n302), .A2(new_n666), .A3(new_n496), .A4(new_n739), .ZN(new_n806));
  INV_X1    g620(.A(new_n420), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n656), .A2(new_n807), .A3(new_n678), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n806), .B(new_n808), .C1(new_n767), .C2(new_n768), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n742), .A2(new_n806), .A3(new_n678), .A4(new_n727), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n769), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n769), .A2(new_n809), .A3(KEYINPUT111), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n577), .B(new_n673), .C1(new_n701), .C2(new_n679), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n760), .A2(new_n666), .A3(new_n700), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n724), .A2(new_n817), .A3(new_n691), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n732), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n816), .A2(new_n732), .A3(new_n821), .A4(new_n818), .ZN(new_n822));
  AND4_X1   g636(.A1(KEYINPUT53), .A2(new_n815), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n744), .A2(new_n758), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n762), .A2(new_n763), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n715), .A2(new_n577), .B1(new_n723), .B2(new_n724), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n709), .A3(new_n712), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n694), .A2(new_n771), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n501), .B(new_n646), .C1(new_n497), .C2(new_n499), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n631), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n503), .B2(new_n667), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT109), .B1(new_n694), .B2(new_n807), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n377), .A2(new_n384), .A3(new_n836), .A4(new_n420), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n832), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n632), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n625), .B(new_n834), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n830), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n828), .A2(new_n709), .A3(new_n712), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n764), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n824), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n823), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n815), .A3(new_n820), .A4(new_n822), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n842), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n852), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n845), .A2(new_n815), .ZN(new_n856));
  INV_X1    g670(.A(new_n842), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n820), .A2(new_n822), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n852), .B1(new_n859), .B2(new_n850), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n853), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n427), .B1(new_n774), .B2(new_n775), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n728), .A2(new_n620), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n708), .A2(new_n502), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT115), .B1(new_n683), .B2(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n683), .A2(KEYINPUT115), .A3(new_n865), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT116), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n706), .A2(new_n301), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT108), .Z(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n707), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n800), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n791), .A3(new_n864), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n759), .A2(new_n189), .A3(new_n872), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n862), .A2(new_n730), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n620), .A2(new_n427), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n692), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n881), .A2(new_n694), .A3(new_n771), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n868), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n871), .A2(new_n877), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n425), .B1(new_n881), .B2(new_n831), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n864), .B2(new_n731), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n862), .A2(new_n757), .A3(new_n878), .ZN(new_n890));
  XOR2_X1   g704(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n891));
  OR2_X1    g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n883), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n871), .A2(new_n896), .A3(new_n886), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n876), .A2(new_n864), .A3(KEYINPUT114), .A4(new_n791), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n864), .A2(new_n791), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n874), .B1(new_n798), .B2(new_n799), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n884), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n895), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n805), .B1(new_n861), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n873), .B(KEYINPUT49), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n637), .A2(new_n189), .A3(new_n502), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n692), .A2(new_n621), .A3(new_n908), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n907), .A2(new_n909), .A3(new_n683), .A4(new_n694), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n804), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n910), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n895), .A2(new_n904), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n859), .A2(new_n850), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT113), .B(new_n854), .C1(new_n914), .C2(new_n852), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n915), .B2(new_n853), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT118), .B(new_n912), .C1(new_n916), .C2(new_n805), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n917), .ZN(G75));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n466), .A2(new_n479), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n477), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n847), .A2(new_n850), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G902), .ZN(new_n924));
  INV_X1    g738(.A(new_n436), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n919), .B(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT119), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n281), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n924), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT56), .B1(new_n930), .B2(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(new_n922), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n927), .A2(new_n932), .ZN(G51));
  NAND2_X1  g747(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n854), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n784), .B(KEYINPUT120), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT57), .Z(new_n937));
  OAI22_X1  g751(.A1(new_n935), .A2(new_n937), .B1(new_n300), .B2(new_n299), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n783), .B(KEYINPUT121), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n928), .B1(new_n938), .B2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  INV_X1    g756(.A(new_n382), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n928), .ZN(G60));
  INV_X1    g760(.A(new_n634), .ZN(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT59), .Z(new_n949));
  AOI211_X1 g763(.A(new_n947), .B(new_n949), .C1(new_n934), .C2(new_n854), .ZN(new_n950));
  INV_X1    g764(.A(new_n949), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n915), .A2(new_n853), .A3(new_n951), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n928), .B(new_n950), .C1(new_n947), .C2(new_n952), .ZN(G63));
  XNOR2_X1  g767(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n847), .B2(new_n850), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(new_n617), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n664), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n929), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G66));
  OAI21_X1  g776(.A(new_n430), .B1(G224), .B2(new_n281), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT123), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n842), .A2(new_n844), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n920), .B1(G898), .B2(new_n281), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  AOI21_X1  g782(.A(new_n802), .B1(new_n779), .B2(new_n793), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n816), .A2(new_n732), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n698), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT62), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n835), .A2(new_n831), .A3(new_n837), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n696), .A2(new_n759), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n974), .C1(new_n622), .C2(new_n624), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n969), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n281), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n546), .B(KEYINPUT124), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n327), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n281), .A2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n827), .A2(new_n769), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT126), .Z(new_n983));
  NAND3_X1  g797(.A1(new_n790), .A2(new_n724), .A3(new_n757), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(new_n969), .A3(new_n970), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n985), .B2(new_n281), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n980), .B1(new_n986), .B2(new_n979), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n986), .B2(new_n979), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n987), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  OAI221_X1 g806(.A(new_n980), .B1(new_n988), .B2(new_n990), .C1(new_n986), .C2(new_n979), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(new_n547), .A2(new_n684), .ZN(new_n995));
  INV_X1    g809(.A(new_n965), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n985), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g811(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n627), .A2(new_n296), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n995), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n976), .A2(new_n996), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n686), .B1(new_n1002), .B2(new_n1000), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n547), .A2(new_n521), .ZN(new_n1004));
  INV_X1    g818(.A(new_n560), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n929), .B1(new_n914), .B2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1001), .A2(new_n1003), .A3(new_n1007), .ZN(G57));
endmodule


